* NGSPICE file created from wrapped_acorn_prng.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

.subckt wrapped_acorn_prng active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ vccd1 vssd1 wb_clk_i
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3155_ _4869_/Q _3074_/A _3153_/Y _3154_/X _3135_/X vssd1 vssd1 vccd1 vccd1 _4869_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3086_ _4861_/Q _3074_/X _3085_/X _3063_/X vssd1 vssd1 vccd1 vccd1 _4861_/D sky130_fd_sc_hd__o211a_1
X_3988_ _4987_/Q _4767_/Q vssd1 vssd1 vccd1 vccd1 _3996_/B sky130_fd_sc_hd__and2_1
X_5216__123 vssd1 vssd1 vccd1 vccd1 _5216__123/HI _5324_/A sky130_fd_sc_hd__conb_1
XFILLER_22_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2939_ _2951_/A _2939_/B vssd1 vssd1 vccd1 vccd1 _2940_/A sky130_fd_sc_hd__and2_1
X_4609_ _4609_/A _4609_/B vssd1 vssd1 vccd1 vccd1 _4610_/A sky130_fd_sc_hd__and2_1
XFILLER_18_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4960_ _4964_/CLK _4960_/D vssd1 vssd1 vccd1 vccd1 _4960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3911_ _3909_/X _3910_/Y _3848_/X vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__a21o_1
X_4891_ _5087_/CLK _4891_/D vssd1 vssd1 vccd1 vccd1 _4891_/Q sky130_fd_sc_hd__dfxtp_1
X_3842_ _3848_/A vssd1 vssd1 vccd1 vccd1 _3842_/X sky130_fd_sc_hd__clkbuf_2
X_3773_ _4076_/A vssd1 vssd1 vccd1 vccd1 _3773_/X sky130_fd_sc_hd__clkbuf_2
X_2724_ _4991_/Q _4783_/Q _2727_/S vssd1 vssd1 vccd1 vccd1 _2725_/B sky130_fd_sc_hd__mux2_1
X_2655_ _2662_/A _2655_/B vssd1 vssd1 vccd1 vccd1 _2656_/A sky130_fd_sc_hd__and2_1
X_4325_ _4325_/A _4325_/B vssd1 vssd1 vccd1 vccd1 _4325_/Y sky130_fd_sc_hd__nand2_1
X_2586_ _2586_/A vssd1 vssd1 vccd1 vccd1 _4743_/D sky130_fd_sc_hd__clkbuf_1
X_4256_ _4284_/A _4256_/B vssd1 vssd1 vccd1 vccd1 _4256_/X sky130_fd_sc_hd__xor2_1
X_3207_ _3233_/A _3207_/B vssd1 vssd1 vccd1 vccd1 _3207_/X sky130_fd_sc_hd__xor2_1
X_4187_ _4281_/A vssd1 vssd1 vccd1 vccd1 _4187_/X sky130_fd_sc_hd__clkbuf_2
X_3138_ _3138_/A _3138_/B _3138_/C vssd1 vssd1 vccd1 vccd1 _3138_/X sky130_fd_sc_hd__and3_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3069_ _4859_/Q _2976_/A _3067_/Y _3068_/X _3037_/X vssd1 vssd1 vccd1 vccd1 _4859_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5177__84 vssd1 vssd1 vccd1 vccd1 _5177__84/HI _5272_/A sky130_fd_sc_hd__conb_1
XFILLER_5_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2440_ _2441_/A vssd1 vssd1 vccd1 vccd1 _2440_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4101_/A _4103_/Y _4108_/X _4052_/A vssd1 vssd1 vccd1 vccd1 _4110_/X sky130_fd_sc_hd__a31o_1
X_5090_ _5091_/CLK _5090_/D vssd1 vssd1 vccd1 vccd1 _5090_/Q sky130_fd_sc_hd__dfxtp_1
X_4041_ _4993_/Q _4773_/Q vssd1 vssd1 vccd1 vccd1 _4042_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _5122_/CLK _4943_/D vssd1 vssd1 vccd1 vccd1 _4943_/Q sky130_fd_sc_hd__dfxtp_1
X_4874_ _5066_/CLK _4874_/D vssd1 vssd1 vccd1 vccd1 _4874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3825_ _4966_/Q _4746_/Q vssd1 vssd1 vccd1 vccd1 _3827_/A sky130_fd_sc_hd__nor2_1
X_3756_ _3753_/X _3754_/Y _3755_/X vssd1 vssd1 vccd1 vccd1 _3756_/X sky130_fd_sc_hd__a21o_1
X_2707_ _2715_/A _2707_/B vssd1 vssd1 vccd1 vccd1 _2708_/A sky130_fd_sc_hd__and2_1
X_3687_ _5114_/Q _4946_/Q _3686_/X _3678_/B vssd1 vssd1 vccd1 vccd1 _3687_/X sky130_fd_sc_hd__a31o_1
X_2638_ _2638_/A vssd1 vssd1 vccd1 vccd1 _4758_/D sky130_fd_sc_hd__clkbuf_1
X_2569_ _2569_/A vssd1 vssd1 vccd1 vccd1 _4738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5288_ _5288_/A _2533_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
X_4308_ _4290_/A _4292_/Y _4297_/B _4305_/A _4295_/Y vssd1 vssd1 vccd1 vccd1 _4308_/Y
+ sky130_fd_sc_hd__a311oi_2
X_4239_ _4239_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4241_/B sky130_fd_sc_hd__and2_1
XFILLER_59_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4590_ _4590_/A vssd1 vssd1 vccd1 vccd1 _5080_/D sky130_fd_sc_hd__clkbuf_1
X_3610_ _4938_/Q _5106_/Q vssd1 vssd1 vccd1 vccd1 _3610_/Y sky130_fd_sc_hd__nand2_1
X_3541_ _3541_/A _3541_/B vssd1 vssd1 vccd1 vccd1 _3546_/A sky130_fd_sc_hd__and2_1
X_3472_ _3466_/A _3466_/B _3471_/Y vssd1 vssd1 vccd1 vccd1 _3477_/A sky130_fd_sc_hd__o21ai_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2423_ _2548_/A vssd1 vssd1 vccd1 vccd1 _2428_/A sky130_fd_sc_hd__buf_6
XFILLER_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5073_ _5098_/CLK _5073_/D vssd1 vssd1 vccd1 vccd1 _5073_/Q sky130_fd_sc_hd__dfxtp_1
X_4024_ _3937_/X _4020_/Y _4021_/X _4023_/X vssd1 vssd1 vccd1 vccd1 _4978_/D sky130_fd_sc_hd__o211a_1
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4926_ _5106_/CLK _4926_/D vssd1 vssd1 vccd1 vccd1 _4926_/Q sky130_fd_sc_hd__dfxtp_1
X_4857_ _5040_/CLK _4857_/D vssd1 vssd1 vccd1 vccd1 _4857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3808_ _3807_/Y _3788_/B _3786_/Y vssd1 vssd1 vccd1 vccd1 _3808_/Y sky130_fd_sc_hd__a21oi_1
X_4788_ _5002_/CLK _4788_/D vssd1 vssd1 vccd1 vccd1 _4788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3739_ _3720_/A _3722_/Y _3728_/B _3736_/A _3726_/Y vssd1 vssd1 vccd1 vccd1 _3739_/Y
+ sky130_fd_sc_hd__a311oi_2
XFILLER_75_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5147__54 vssd1 vssd1 vccd1 vccd1 _5147__54/HI _5242_/A sky130_fd_sc_hd__conb_1
XFILLER_3_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2972_ _3168_/A _4844_/Q _4845_/Q vssd1 vssd1 vccd1 vccd1 _4129_/A sky130_fd_sc_hd__or3b_4
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4711_ _4711_/A vssd1 vssd1 vccd1 vccd1 _5115_/D sky130_fd_sc_hd__clkbuf_1
X_4642_ _4642_/A vssd1 vssd1 vccd1 vccd1 _5095_/D sky130_fd_sc_hd__clkbuf_1
X_4573_ _4573_/A vssd1 vssd1 vccd1 vccd1 _5075_/D sky130_fd_sc_hd__clkbuf_1
X_3524_ _3523_/Y _3499_/Y _3522_/B _3500_/A vssd1 vssd1 vccd1 vccd1 _3524_/Y sky130_fd_sc_hd__a211oi_1
X_3455_ _4219_/A _3553_/B vssd1 vssd1 vccd1 vccd1 _3544_/B sky130_fd_sc_hd__nor2_2
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3386_ _4911_/Q _5079_/Q vssd1 vssd1 vccd1 vccd1 _3388_/A sky130_fd_sc_hd__nor2_1
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5056_ _5058_/CLK _5056_/D vssd1 vssd1 vccd1 vccd1 _5056_/Q sky130_fd_sc_hd__dfxtp_1
X_4007_ _4976_/Q _3933_/X _4006_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _4976_/D sky130_fd_sc_hd__o211a_1
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4909_ _5091_/CLK _4909_/D vssd1 vssd1 vccd1 vccd1 _4909_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_14_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5018_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _4892_/Q _5060_/Q vssd1 vssd1 vccd1 vccd1 _3241_/B sky130_fd_sc_hd__or2_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3257_/B vssd1 vssd1 vccd1 vccd1 _3223_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2955_ _4418_/A _2955_/B vssd1 vssd1 vccd1 vccd1 _2956_/A sky130_fd_sc_hd__and2_1
X_2886_ _2889_/A vssd1 vssd1 vccd1 vccd1 _2886_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4625_ _4911_/Q _5091_/Q _4629_/S vssd1 vssd1 vccd1 vccd1 _4626_/B sky130_fd_sc_hd__mux2_1
X_4556_ _4891_/Q _5071_/Q _4561_/S vssd1 vssd1 vccd1 vccd1 _4557_/B sky130_fd_sc_hd__mux2_1
X_3507_ _3521_/A _3508_/B vssd1 vssd1 vccd1 vccd1 _3507_/X sky130_fd_sc_hd__or2_1
X_4487_ _4871_/Q _5051_/Q _4491_/S vssd1 vssd1 vccd1 vccd1 _4488_/B sky130_fd_sc_hd__mux2_1
X_3438_ _3436_/Y _3438_/B vssd1 vssd1 vccd1 vccd1 _3438_/X sky130_fd_sc_hd__and2b_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _4896_/Q _3363_/X _3368_/X _3353_/X vssd1 vssd1 vccd1 vccd1 _4896_/D sky130_fd_sc_hd__o211a_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5121_/CLK _5108_/D vssd1 vssd1 vccd1 vccd1 _5108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5039_ _5040_/CLK _5039_/D vssd1 vssd1 vccd1 vccd1 _5039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2740_ _2750_/A _2740_/B vssd1 vssd1 vccd1 vccd1 _2741_/A sky130_fd_sc_hd__and2_1
X_2671_ _4976_/Q _4768_/Q _2674_/S vssd1 vssd1 vccd1 vccd1 _2672_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4410_ _4410_/A vssd1 vssd1 vccd1 vccd1 _5028_/D sky130_fd_sc_hd__clkbuf_1
X_4341_ _4341_/A _4341_/B vssd1 vssd1 vccd1 vccd1 _4341_/Y sky130_fd_sc_hd__nor2_1
X_4272_ _4271_/Y _4263_/B _4269_/Y vssd1 vssd1 vccd1 vccd1 _4272_/Y sky130_fd_sc_hd__a21oi_1
X_3223_ _3223_/A _3223_/B vssd1 vssd1 vccd1 vccd1 _3223_/Y sky130_fd_sc_hd__nand2_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3154_ _3144_/A _3146_/Y _3152_/X _3084_/A vssd1 vssd1 vccd1 vccd1 _3154_/X sky130_fd_sc_hd__a31o_1
X_3085_ _3082_/X _3083_/Y _3084_/X vssd1 vssd1 vccd1 vccd1 _3085_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3987_ _4986_/Q _4766_/Q vssd1 vssd1 vccd1 vccd1 _3995_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2938_ _5279_/A _4854_/Q _2944_/S vssd1 vssd1 vccd1 vccd1 _2939_/B sky130_fd_sc_hd__mux2_1
X_2869_ _3037_/A vssd1 vssd1 vccd1 vccd1 _2869_/X sky130_fd_sc_hd__clkbuf_2
X_4608_ _4906_/Q _5086_/Q _4612_/S vssd1 vssd1 vccd1 vccd1 _4609_/B sky130_fd_sc_hd__mux2_1
X_4539_ _4539_/A _4539_/B vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__and2_1
XFILLER_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5198__105 vssd1 vssd1 vccd1 vccd1 _5198__105/HI _5306_/A sky130_fd_sc_hd__conb_1
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3910_ _3910_/A _3910_/B vssd1 vssd1 vccd1 vccd1 _3910_/Y sky130_fd_sc_hd__nand2_2
X_4890_ _5070_/CLK _4890_/D vssd1 vssd1 vccd1 vccd1 _4890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3841_ _4219_/A _3936_/B vssd1 vssd1 vccd1 vccd1 _3848_/A sky130_fd_sc_hd__or2_2
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3772_ _3763_/A _3765_/Y _3770_/Y _3755_/X vssd1 vssd1 vccd1 vccd1 _3772_/X sky130_fd_sc_hd__a31o_1
X_2723_ _2723_/A vssd1 vssd1 vccd1 vccd1 _4782_/D sky130_fd_sc_hd__clkbuf_1
X_2654_ _4971_/Q _4763_/Q _2657_/S vssd1 vssd1 vccd1 vccd1 _2655_/B sky130_fd_sc_hd__mux2_1
X_2585_ _2592_/A _2585_/B vssd1 vssd1 vccd1 vccd1 _2586_/A sky130_fd_sc_hd__and2_1
X_4324_ _4325_/A _4325_/B vssd1 vssd1 vccd1 vccd1 _4324_/X sky130_fd_sc_hd__or2_1
XFILLER_59_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4255_ _4241_/A _4241_/B _4246_/Y _4254_/X vssd1 vssd1 vccd1 vccd1 _4256_/B sky130_fd_sc_hd__a31o_1
X_4186_ _4182_/Y _4176_/X _4189_/B _4191_/C _4136_/A vssd1 vssd1 vccd1 vccd1 _4186_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_67_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3206_ _3191_/A _3191_/B _3197_/Y _3205_/X vssd1 vssd1 vccd1 vccd1 _3207_/B sky130_fd_sc_hd__a31o_1
X_3137_ _3137_/A _3137_/B _3139_/C vssd1 vssd1 vccd1 vccd1 _3138_/C sky130_fd_sc_hd__and3_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3068_ _3059_/B _3065_/X _3066_/X _2988_/A vssd1 vssd1 vccd1 vccd1 _3068_/X sky130_fd_sc_hd__a31o_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5192__99 vssd1 vssd1 vccd1 vccd1 _5192__99/HI _5300_/A sky130_fd_sc_hd__conb_1
XFILLER_78_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4040_ _4980_/Q _4034_/X _4039_/X _4023_/X vssd1 vssd1 vccd1 vccd1 _4980_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4942_ _5121_/CLK _4942_/D vssd1 vssd1 vccd1 vccd1 _4942_/Q sky130_fd_sc_hd__dfxtp_1
X_4873_ _5066_/CLK _4873_/D vssd1 vssd1 vccd1 vccd1 _4873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3824_ _4953_/Q _3784_/X _3822_/Y _3823_/X _3773_/X vssd1 vssd1 vccd1 vccd1 _4953_/D
+ sky130_fd_sc_hd__o221a_1
X_3755_ _3755_/A vssd1 vssd1 vccd1 vccd1 _3755_/X sky130_fd_sc_hd__clkbuf_2
X_2706_ _4986_/Q _4778_/Q _2710_/S vssd1 vssd1 vccd1 vccd1 _2707_/B sky130_fd_sc_hd__mux2_1
X_3686_ _5115_/Q _4947_/Q vssd1 vssd1 vccd1 vccd1 _3686_/X sky130_fd_sc_hd__or2_1
X_2637_ _2645_/A _2637_/B vssd1 vssd1 vccd1 vccd1 _2638_/A sky130_fd_sc_hd__and2_1
X_2568_ _2575_/A _2568_/B vssd1 vssd1 vccd1 vccd1 _2569_/A sky130_fd_sc_hd__and2_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5287_ _5287_/A _2483_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
X_2499_ _2503_/A vssd1 vssd1 vccd1 vccd1 _2499_/Y sky130_fd_sc_hd__inv_2
X_4307_ _4224_/X _4305_/X _4306_/X _4232_/X vssd1 vssd1 vccd1 vccd1 _5014_/D sky130_fd_sc_hd__o211a_1
X_4238_ _5018_/Q _4798_/Q vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__or2_1
X_4169_ _4169_/A _4169_/B vssd1 vssd1 vccd1 vccd1 _4190_/B sky130_fd_sc_hd__and2_1
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5098_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3540_ _4930_/Q _5098_/Q vssd1 vssd1 vccd1 vccd1 _3541_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3471_ _4921_/Q _5089_/Q vssd1 vssd1 vccd1 vccd1 _3471_/Y sky130_fd_sc_hd__nand2_1
X_2422_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2422_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5072_ _5087_/CLK _5072_/D vssd1 vssd1 vccd1 vccd1 _5072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4023_ _4321_/A vssd1 vssd1 vccd1 vccd1 _4023_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4925_ _5106_/CLK _4925_/D vssd1 vssd1 vccd1 vccd1 _4925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4856_ _5041_/CLK _4856_/D vssd1 vssd1 vccd1 vccd1 _4856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3807_ _4960_/Q _4740_/Q vssd1 vssd1 vccd1 vccd1 _3807_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4787_ _5002_/CLK _4787_/D vssd1 vssd1 vccd1 vccd1 _4787_/Q sky130_fd_sc_hd__dfxtp_1
X_3738_ _3656_/X _3736_/X _3737_/X _3724_/X vssd1 vssd1 vccd1 vccd1 _4942_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3669_ _5114_/Q _4946_/Q vssd1 vssd1 vccd1 vccd1 _3671_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5162__69 vssd1 vssd1 vccd1 vccd1 _5162__69/HI _5257_/A sky130_fd_sc_hd__conb_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2971_ _3077_/B vssd1 vssd1 vccd1 vccd1 _3175_/A sky130_fd_sc_hd__clkbuf_2
X_4710_ _4713_/A _4710_/B vssd1 vssd1 vccd1 vccd1 _4711_/A sky130_fd_sc_hd__and2_1
X_4641_ _4644_/A _4641_/B vssd1 vssd1 vccd1 vccd1 _4642_/A sky130_fd_sc_hd__and2_1
X_4572_ _4575_/A _4572_/B vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__and2_1
X_3523_ _4924_/Q _5092_/Q vssd1 vssd1 vccd1 vccd1 _3523_/Y sky130_fd_sc_hd__nand2_1
X_3454_ _4907_/Q _3401_/X _3452_/X _3453_/Y _3441_/X vssd1 vssd1 vccd1 vccd1 _4907_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3385_ _3376_/Y _3367_/X _3384_/Y _2967_/A vssd1 vssd1 vccd1 vccd1 _4898_/D sky130_fd_sc_hd__a211oi_1
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5055_ _5066_/CLK _5055_/D vssd1 vssd1 vccd1 vccd1 _5055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4006_ _4004_/Y _4005_/X _3943_/X vssd1 vssd1 vccd1 vccd1 _4006_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4908_ _5091_/CLK _4908_/D vssd1 vssd1 vccd1 vccd1 _4908_/Q sky130_fd_sc_hd__dfxtp_1
X_4839_ _5033_/CLK _4839_/D vssd1 vssd1 vccd1 vccd1 _5280_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3175_/A _4318_/A vssd1 vssd1 vccd1 vccd1 _3257_/B sky130_fd_sc_hd__nor2_2
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2954_ _5284_/A _4859_/Q _2954_/S vssd1 vssd1 vccd1 vccd1 _2955_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2885_ _2878_/X _4825_/Q _2882_/X _2884_/X _2876_/X vssd1 vssd1 vccd1 vccd1 _4825_/D
+ sky130_fd_sc_hd__o221a_1
X_4624_ _4624_/A vssd1 vssd1 vccd1 vccd1 _5090_/D sky130_fd_sc_hd__clkbuf_1
X_4555_ _4555_/A vssd1 vssd1 vccd1 vccd1 _5070_/D sky130_fd_sc_hd__clkbuf_1
X_3506_ _3501_/A _3499_/Y _3500_/A vssd1 vssd1 vccd1 vccd1 _3508_/B sky130_fd_sc_hd__a21o_1
X_4486_ _4486_/A vssd1 vssd1 vccd1 vccd1 _5050_/D sky130_fd_sc_hd__clkbuf_1
X_3437_ _4917_/Q _5085_/Q vssd1 vssd1 vccd1 vccd1 _3438_/B sky130_fd_sc_hd__nand2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3364_/X _3372_/A _3367_/X vssd1 vssd1 vccd1 vccd1 _3368_/X sky130_fd_sc_hd__a21o_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5107_ _5107_/CLK _5107_/D vssd1 vssd1 vccd1 vccd1 _5107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3299_ _3299_/A _3299_/B vssd1 vssd1 vccd1 vccd1 _3328_/A sky130_fd_sc_hd__nor2_1
X_5038_ _5040_/CLK _5038_/D vssd1 vssd1 vccd1 vccd1 _5038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5132__39 vssd1 vssd1 vccd1 vccd1 _5132__39/HI _5227_/A sky130_fd_sc_hd__conb_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5200__107 vssd1 vssd1 vccd1 vccd1 _5200__107/HI _5308_/A sky130_fd_sc_hd__conb_1
XFILLER_29_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2670_ _2670_/A vssd1 vssd1 vccd1 vccd1 _4767_/D sky130_fd_sc_hd__clkbuf_1
X_4340_ _4823_/Q _4811_/Q vssd1 vssd1 vccd1 vccd1 _4341_/B sky130_fd_sc_hd__and2_1
X_4271_ _5020_/Q _4800_/Q vssd1 vssd1 vccd1 vccd1 _4271_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3222_ _3225_/A _3225_/B vssd1 vssd1 vccd1 vccd1 _3223_/B sky130_fd_sc_hd__xnor2_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3153_ _3144_/A _3146_/Y _3152_/X vssd1 vssd1 vccd1 vccd1 _3153_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3084_ _3084_/A vssd1 vssd1 vccd1 vccd1 _3084_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3986_ _4974_/Q _3933_/X _3985_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _4974_/D sky130_fd_sc_hd__o211a_1
X_2937_ _4454_/A vssd1 vssd1 vccd1 vccd1 _2951_/A sky130_fd_sc_hd__clkbuf_2
X_4607_ _4607_/A vssd1 vssd1 vccd1 vccd1 _5085_/D sky130_fd_sc_hd__clkbuf_1
X_2868_ _2982_/A vssd1 vssd1 vccd1 vccd1 _3037_/A sky130_fd_sc_hd__clkbuf_2
X_2799_ _2803_/A _2799_/B vssd1 vssd1 vccd1 vccd1 _2800_/A sky130_fd_sc_hd__and2_1
X_4538_ _4886_/Q _5066_/Q _4542_/S vssd1 vssd1 vccd1 vccd1 _4539_/B sky130_fd_sc_hd__mux2_1
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4469_ _4866_/Q _5046_/Q _4474_/S vssd1 vssd1 vccd1 vccd1 _4470_/B sky130_fd_sc_hd__mux2_1
XFILLER_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ _4968_/Q _4748_/Q vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3771_ _3763_/A _3765_/Y _3770_/Y vssd1 vssd1 vccd1 vccd1 _3771_/Y sky130_fd_sc_hd__a21oi_1
X_2722_ _2733_/A _2722_/B vssd1 vssd1 vccd1 vccd1 _2723_/A sky130_fd_sc_hd__and2_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2653_ _2653_/A vssd1 vssd1 vccd1 vccd1 _4762_/D sky130_fd_sc_hd__clkbuf_1
X_2584_ _4951_/Q _4743_/Q _2587_/S vssd1 vssd1 vccd1 vccd1 _2585_/B sky130_fd_sc_hd__mux2_1
X_4323_ _4821_/Q _4809_/Q vssd1 vssd1 vccd1 vccd1 _4325_/B sky130_fd_sc_hd__xnor2_1
X_4254_ _5018_/Q _4798_/Q _4253_/X _4246_/B vssd1 vssd1 vccd1 vccd1 _4254_/X sky130_fd_sc_hd__a31o_1
X_4185_ _4182_/Y _4176_/X _4189_/B _4191_/C vssd1 vssd1 vccd1 vccd1 _4185_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3205_ _4886_/Q _5054_/Q _3204_/X _3197_/B vssd1 vssd1 vccd1 vccd1 _3205_/X sky130_fd_sc_hd__a31o_1
XFILLER_67_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3136_ _4867_/Q _3074_/A _3131_/Y _3132_/X _3135_/X vssd1 vssd1 vccd1 vccd1 _4867_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3067_ _3059_/B _3065_/X _3066_/X vssd1 vssd1 vccd1 vccd1 _3067_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3969_ _3954_/A _3954_/B _3959_/Y _3968_/X vssd1 vssd1 vccd1 vccd1 _3971_/B sky130_fd_sc_hd__a31o_1
XFILLER_5_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5206__113 vssd1 vssd1 vccd1 vccd1 _5206__113/HI _5314_/A sky130_fd_sc_hd__conb_1
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4941_ _5121_/CLK _4941_/D vssd1 vssd1 vccd1 vccd1 _4941_/Q sky130_fd_sc_hd__dfxtp_1
X_4872_ _5048_/CLK _4872_/D vssd1 vssd1 vccd1 vccd1 _4872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3823_ _3814_/A _3816_/Y _3821_/X _3755_/A vssd1 vssd1 vccd1 vccd1 _3823_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5002_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3754_ _3754_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _3754_/Y sky130_fd_sc_hd__nand2_1
X_2705_ _2705_/A vssd1 vssd1 vccd1 vccd1 _4777_/D sky130_fd_sc_hd__clkbuf_1
X_5168__75 vssd1 vssd1 vccd1 vccd1 _5168__75/HI _5263_/A sky130_fd_sc_hd__conb_1
X_3685_ _3685_/A _3685_/B vssd1 vssd1 vccd1 vccd1 _3712_/A sky130_fd_sc_hd__nor2_1
X_2636_ _4966_/Q _4758_/Q _2639_/S vssd1 vssd1 vccd1 vccd1 _2637_/B sky130_fd_sc_hd__mux2_1
X_2567_ _4946_/Q _4738_/Q _2570_/S vssd1 vssd1 vccd1 vccd1 _2568_/B sky130_fd_sc_hd__mux2_1
X_5286_ _5286_/A _2482_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
X_2498_ _2516_/A vssd1 vssd1 vccd1 vccd1 _2503_/A sky130_fd_sc_hd__buf_8
X_4306_ _5014_/Q _4306_/B vssd1 vssd1 vccd1 vccd1 _4306_/X sky130_fd_sc_hd__or2_1
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4237_ _5018_/Q _4798_/Q vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__nand2_1
XFILLER_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4168_ _5009_/Q _4789_/Q vssd1 vssd1 vccd1 vccd1 _4169_/B sky130_fd_sc_hd__nand2_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4099_ _5000_/Q _4780_/Q vssd1 vssd1 vccd1 vccd1 _4101_/A sky130_fd_sc_hd__nand2_1
X_3119_ _4878_/Q _5046_/Q vssd1 vssd1 vccd1 vccd1 _3137_/A sky130_fd_sc_hd__xor2_1
XFILLER_55_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3470_ _4910_/Q vssd1 vssd1 vccd1 vccd1 _3470_/Y sky130_fd_sc_hd__inv_2
X_2421_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2421_/Y sky130_fd_sc_hd__inv_2
X_5071_ _5085_/CLK _5071_/D vssd1 vssd1 vccd1 vccd1 _5071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4022_ _4022_/A vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__buf_2
XFILLER_37_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4924_ _5106_/CLK _4924_/D vssd1 vssd1 vccd1 vccd1 _4924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4855_ _5046_/CLK _4855_/D vssd1 vssd1 vccd1 vccd1 _4855_/Q sky130_fd_sc_hd__dfxtp_1
X_4786_ _4995_/CLK _4786_/D vssd1 vssd1 vccd1 vccd1 _4786_/Q sky130_fd_sc_hd__dfxtp_1
X_3806_ _3806_/A _3806_/B _3806_/C vssd1 vssd1 vccd1 vccd1 _3806_/X sky130_fd_sc_hd__and3_1
X_3737_ _4942_/Q _3737_/B vssd1 vssd1 vccd1 vccd1 _3737_/X sky130_fd_sc_hd__or2_1
X_3668_ _3663_/A _3663_/B _3667_/Y vssd1 vssd1 vccd1 vccd1 _3673_/A sky130_fd_sc_hd__o21ai_1
X_2619_ _4961_/Q _4753_/Q _2622_/S vssd1 vssd1 vccd1 vccd1 _2620_/B sky130_fd_sc_hd__mux2_1
X_3599_ _3598_/A _3617_/B _3564_/X vssd1 vssd1 vccd1 vccd1 _3599_/X sky130_fd_sc_hd__a21o_1
X_5269_ _5269_/A _2462_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2970_ _3648_/A _4030_/B vssd1 vssd1 vccd1 vccd1 _3077_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _4915_/Q _5095_/Q _4648_/S vssd1 vssd1 vccd1 vccd1 _4641_/B sky130_fd_sc_hd__mux2_1
X_4571_ _4895_/Q _5075_/Q _4578_/S vssd1 vssd1 vccd1 vccd1 _4572_/B sky130_fd_sc_hd__mux2_1
X_5138__45 vssd1 vssd1 vccd1 vccd1 _5138__45/HI _5233_/A sky130_fd_sc_hd__conb_1
X_3522_ _3522_/A _3522_/B vssd1 vssd1 vccd1 vccd1 _3522_/Y sky130_fd_sc_hd__nor2_1
X_3453_ _3445_/B _3450_/Y _3451_/Y _3401_/X vssd1 vssd1 vccd1 vccd1 _3453_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3384_ _3382_/X _3383_/Y _3367_/X vssd1 vssd1 vccd1 vccd1 _3384_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5066_/CLK _5054_/D vssd1 vssd1 vccd1 vccd1 _5054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4005_ _4004_/A _4004_/B _4004_/C vssd1 vssd1 vccd1 vccd1 _4005_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4907_ _5098_/CLK _4907_/D vssd1 vssd1 vccd1 vccd1 _4907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4838_ _5033_/CLK _4838_/D vssd1 vssd1 vccd1 vccd1 _5279_/A sky130_fd_sc_hd__dfxtp_1
X_4769_ _4975_/CLK _4769_/D vssd1 vssd1 vccd1 vccd1 _4769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4948_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2953_ _4454_/A vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__buf_2
X_2884_ _2865_/X input23/X _2883_/X vssd1 vssd1 vccd1 vccd1 _2884_/X sky130_fd_sc_hd__a21bo_1
X_4623_ _4626_/A _4623_/B vssd1 vssd1 vccd1 vccd1 _4624_/A sky130_fd_sc_hd__and2_1
X_4554_ _4557_/A _4554_/B vssd1 vssd1 vccd1 vccd1 _4555_/A sky130_fd_sc_hd__and2_1
X_3505_ _4926_/Q _5094_/Q vssd1 vssd1 vccd1 vccd1 _3521_/A sky130_fd_sc_hd__xnor2_1
X_4485_ _4488_/A _4485_/B vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__and2_1
X_3436_ _4917_/Q _5085_/Q vssd1 vssd1 vccd1 vccd1 _3436_/Y sky130_fd_sc_hd__nor2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3373_/A vssd1 vssd1 vccd1 vccd1 _3367_/X sky130_fd_sc_hd__clkbuf_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5106_/CLK _5106_/D vssd1 vssd1 vccd1 vccd1 _5106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3298_ _4900_/Q _5068_/Q vssd1 vssd1 vccd1 vccd1 _3299_/B sky130_fd_sc_hd__nor2_1
X_5037_ _5040_/CLK _5037_/D vssd1 vssd1 vccd1 vccd1 _5037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4270_ _4264_/A _4263_/B _4268_/Y _4269_/Y vssd1 vssd1 vccd1 vccd1 _4270_/X sky130_fd_sc_hd__a211o_1
X_3221_ _3215_/A _3214_/B _3212_/Y vssd1 vssd1 vccd1 vccd1 _3225_/B sky130_fd_sc_hd__a21o_1
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3152_ _3150_/Y _3152_/B vssd1 vssd1 vccd1 vccd1 _3152_/X sky130_fd_sc_hd__and2b_1
X_3083_ _3083_/A _3083_/B vssd1 vssd1 vccd1 vccd1 _3083_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3985_ _3983_/X _3984_/Y _3943_/X vssd1 vssd1 vccd1 vccd1 _3985_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2936_ _4646_/A vssd1 vssd1 vccd1 vccd1 _4454_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2867_ _2865_/X input19/X _2878_/A vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__a21bo_1
X_4606_ _4609_/A _4606_/B vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__and2_1
X_2798_ _5012_/Q _4804_/Q _2798_/S vssd1 vssd1 vccd1 vccd1 _2799_/B sky130_fd_sc_hd__mux2_1
X_4537_ _4537_/A vssd1 vssd1 vccd1 vccd1 _5065_/D sky130_fd_sc_hd__clkbuf_1
X_4468_ _4468_/A vssd1 vssd1 vccd1 vccd1 _5045_/D sky130_fd_sc_hd__clkbuf_1
X_3419_ _3421_/B _3421_/C _3417_/Y _3373_/A vssd1 vssd1 vccd1 vccd1 _3419_/X sky130_fd_sc_hd__a31o_1
X_4399_ _4399_/A _4399_/B vssd1 vssd1 vccd1 vccd1 _4399_/X sky130_fd_sc_hd__xor2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3770_ _3770_/A _3770_/B vssd1 vssd1 vccd1 vccd1 _3770_/Y sky130_fd_sc_hd__nor2_1
X_2721_ _4990_/Q _4782_/Q _2727_/S vssd1 vssd1 vccd1 vccd1 _2722_/B sky130_fd_sc_hd__mux2_1
XFILLER_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2652_ _2662_/A _2652_/B vssd1 vssd1 vccd1 vccd1 _2653_/A sky130_fd_sc_hd__and2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2583_ _2583_/A vssd1 vssd1 vccd1 vccd1 _4742_/D sky130_fd_sc_hd__clkbuf_1
X_4322_ _5016_/Q _4315_/X _4320_/X _4321_/X vssd1 vssd1 vccd1 vccd1 _5016_/D sky130_fd_sc_hd__o211a_1
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4253_ _5019_/Q _4799_/Q vssd1 vssd1 vccd1 vccd1 _4253_/X sky130_fd_sc_hd__or2_1
X_3204_ _4887_/Q _5055_/Q vssd1 vssd1 vccd1 vccd1 _3204_/X sky130_fd_sc_hd__or2_1
X_4184_ _5011_/Q _4791_/Q vssd1 vssd1 vccd1 vccd1 _4191_/C sky130_fd_sc_hd__or2_1
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3135_ _3551_/A vssd1 vssd1 vccd1 vccd1 _3135_/X sky130_fd_sc_hd__buf_2
XFILLER_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3066_ _4871_/Q _5039_/Q vssd1 vssd1 vccd1 vccd1 _3066_/X sky130_fd_sc_hd__xor2_1
XFILLER_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3968_ _4982_/Q _4762_/Q _3967_/X _3959_/B vssd1 vssd1 vccd1 vccd1 _3968_/X sky130_fd_sc_hd__a31o_1
XFILLER_23_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2919_ _2919_/A vssd1 vssd1 vccd1 vccd1 _2934_/A sky130_fd_sc_hd__clkbuf_2
X_3899_ _3895_/Y _3889_/X _3901_/B _3903_/C _3848_/A vssd1 vssd1 vccd1 vccd1 _3899_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4940_ _5121_/CLK _4940_/D vssd1 vssd1 vccd1 vccd1 _4940_/Q sky130_fd_sc_hd__dfxtp_1
X_4871_ _5050_/CLK _4871_/D vssd1 vssd1 vccd1 vccd1 _4871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3822_ _3814_/A _3816_/Y _3821_/X vssd1 vssd1 vccd1 vccd1 _3822_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3753_ _3754_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _3753_/X sky130_fd_sc_hd__or2_1
X_2704_ _2715_/A _2704_/B vssd1 vssd1 vccd1 vccd1 _2705_/A sky130_fd_sc_hd__and2_1
X_3684_ _5116_/Q _4948_/Q vssd1 vssd1 vccd1 vccd1 _3685_/B sky130_fd_sc_hd__nor2_1
X_2635_ _2635_/A vssd1 vssd1 vccd1 vccd1 _4757_/D sky130_fd_sc_hd__clkbuf_1
X_4305_ _4305_/A _4305_/B vssd1 vssd1 vccd1 vccd1 _4305_/X sky130_fd_sc_hd__xor2_1
X_2566_ _2566_/A vssd1 vssd1 vccd1 vccd1 _4737_/D sky130_fd_sc_hd__clkbuf_1
X_5285_ _5285_/A _2481_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
X_2497_ _2497_/A vssd1 vssd1 vccd1 vccd1 _2497_/Y sky130_fd_sc_hd__inv_2
X_4236_ _4229_/A _4229_/B _4235_/Y vssd1 vssd1 vccd1 vccd1 _4241_/A sky130_fd_sc_hd__o21ai_1
X_4167_ _5009_/Q _4789_/Q vssd1 vssd1 vccd1 vccd1 _4169_/A sky130_fd_sc_hd__or2_1
X_3118_ _4865_/Q _3074_/A _3116_/Y _3117_/X _3037_/X vssd1 vssd1 vccd1 vccd1 _4865_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_55_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4098_ _4067_/B _4093_/X _4097_/X vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__a21o_1
XFILLER_70_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3049_ _3047_/X _3048_/Y _2988_/X vssd1 vssd1 vccd1 vccd1 _3049_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_48_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5032_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2420_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2420_/Y sky130_fd_sc_hd__inv_2
X_5070_ _5070_/CLK _5070_/D vssd1 vssd1 vccd1 vccd1 _5070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4021_ _4978_/Q _4021_/B vssd1 vssd1 vccd1 vccd1 _4021_/X sky130_fd_sc_hd__or2_1
XFILLER_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4923_ _5106_/CLK _4923_/D vssd1 vssd1 vccd1 vccd1 _4923_/Q sky130_fd_sc_hd__dfxtp_1
X_4854_ _5041_/CLK _4854_/D vssd1 vssd1 vccd1 vccd1 _4854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4785_ _5002_/CLK _4785_/D vssd1 vssd1 vccd1 vccd1 _4785_/Q sky130_fd_sc_hd__dfxtp_1
X_3805_ _3805_/A _3805_/B _3805_/C vssd1 vssd1 vccd1 vccd1 _3806_/C sky130_fd_sc_hd__and3_1
X_3736_ _3736_/A _3736_/B vssd1 vssd1 vccd1 vccd1 _3736_/X sky130_fd_sc_hd__xor2_1
X_3667_ _5113_/Q _4945_/Q vssd1 vssd1 vccd1 vccd1 _3667_/Y sky130_fd_sc_hd__nand2_1
X_2618_ _2618_/A vssd1 vssd1 vccd1 vccd1 _4752_/D sky130_fd_sc_hd__clkbuf_1
X_3598_ _3598_/A _3617_/B vssd1 vssd1 vccd1 vccd1 _3598_/Y sky130_fd_sc_hd__nor2_1
X_2549_ _5285_/A vssd1 vssd1 vccd1 vccd1 _3133_/A sky130_fd_sc_hd__inv_2
X_5268_ _5268_/A _2459_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
X_4219_ _4219_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _4306_/B sky130_fd_sc_hd__nor2_2
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4570_ _4570_/A vssd1 vssd1 vccd1 vccd1 _5074_/D sky130_fd_sc_hd__clkbuf_1
X_3521_ _3521_/A _3521_/B _3521_/C vssd1 vssd1 vccd1 vccd1 _3522_/B sky130_fd_sc_hd__or3_1
X_3452_ _3445_/B _3450_/Y _3451_/Y vssd1 vssd1 vccd1 vccd1 _3452_/X sky130_fd_sc_hd__o21a_1
X_3383_ _3383_/A _3383_/B vssd1 vssd1 vccd1 vccd1 _3383_/Y sky130_fd_sc_hd__nand2_1
X_5122_ _5122_/CLK _5122_/D vssd1 vssd1 vccd1 vccd1 _5122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5053_ _5066_/CLK _5053_/D vssd1 vssd1 vccd1 vccd1 _5053_/Q sky130_fd_sc_hd__dfxtp_1
X_4004_ _4004_/A _4004_/B _4004_/C vssd1 vssd1 vccd1 vccd1 _4004_/Y sky130_fd_sc_hd__nand3_1
XFILLER_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _5085_/CLK _4906_/D vssd1 vssd1 vccd1 vccd1 _4906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4837_ _5033_/CLK _4837_/D vssd1 vssd1 vccd1 vccd1 _5278_/A sky130_fd_sc_hd__dfxtp_1
X_4768_ _4975_/CLK _4768_/D vssd1 vssd1 vccd1 vccd1 _4768_/Q sky130_fd_sc_hd__dfxtp_1
X_4699_ _4932_/Q _5112_/Q _4699_/S vssd1 vssd1 vccd1 vccd1 _4700_/B sky130_fd_sc_hd__mux2_1
X_3719_ _5120_/Q _4952_/Q vssd1 vssd1 vccd1 vccd1 _3720_/B sky130_fd_sc_hd__or2_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2952_ _2952_/A vssd1 vssd1 vccd1 vccd1 _4842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2883_ _2958_/B vssd1 vssd1 vccd1 vccd1 _2883_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4622_ _4910_/Q _5090_/Q _4629_/S vssd1 vssd1 vccd1 vccd1 _4623_/B sky130_fd_sc_hd__mux2_1
X_4553_ _4890_/Q _5070_/Q _4561_/S vssd1 vssd1 vccd1 vccd1 _4554_/B sky130_fd_sc_hd__mux2_1
X_3504_ _3461_/X _3501_/X _3502_/X _3503_/X vssd1 vssd1 vccd1 vccd1 _4913_/D sky130_fd_sc_hd__o211a_1
X_4484_ _4870_/Q _5050_/Q _4491_/S vssd1 vssd1 vccd1 vccd1 _4485_/B sky130_fd_sc_hd__mux2_1
X_3435_ _4904_/Q _3363_/X _3433_/X _3434_/X vssd1 vssd1 vccd1 vccd1 _4904_/D sky130_fd_sc_hd__o211a_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _4125_/A _3557_/B vssd1 vssd1 vccd1 vccd1 _3373_/A sky130_fd_sc_hd__or2_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _4900_/Q _5068_/Q vssd1 vssd1 vccd1 vccd1 _3299_/A sky130_fd_sc_hd__and2_1
X_5105_ _5106_/CLK _5105_/D vssd1 vssd1 vccd1 vccd1 _5105_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5041_/CLK _5036_/D vssd1 vssd1 vccd1 vccd1 _5036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3220_ _3232_/A _3232_/B vssd1 vssd1 vccd1 vccd1 _3225_/A sky130_fd_sc_hd__nand2_1
XFILLER_79_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3151_ _4881_/Q _5049_/Q vssd1 vssd1 vccd1 vccd1 _3152_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3082_ _3083_/A _3083_/B vssd1 vssd1 vccd1 vccd1 _3082_/X sky130_fd_sc_hd__or2_1
XFILLER_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3984_ _3996_/A _3984_/B vssd1 vssd1 vccd1 vccd1 _3984_/Y sky130_fd_sc_hd__nand2_1
X_2935_ _2935_/A vssd1 vssd1 vccd1 vccd1 _4837_/D sky130_fd_sc_hd__clkbuf_1
X_2866_ _2958_/B vssd1 vssd1 vccd1 vccd1 _2878_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4605_ _4905_/Q _5085_/Q _4612_/S vssd1 vssd1 vccd1 vccd1 _4606_/B sky130_fd_sc_hd__mux2_1
XFILLER_7_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2797_ _2797_/A vssd1 vssd1 vccd1 vccd1 _4803_/D sky130_fd_sc_hd__clkbuf_1
X_4536_ _4539_/A _4536_/B vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__and2_1
X_4467_ _4470_/A _4467_/B vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__and2_1
X_3418_ _3421_/B _3421_/C _3417_/Y vssd1 vssd1 vccd1 vccd1 _3418_/Y sky130_fd_sc_hd__a21oi_1
X_4398_ _4384_/A _4386_/Y _4391_/B _4389_/Y vssd1 vssd1 vccd1 vccd1 _4399_/B sky130_fd_sc_hd__a31o_1
X_3349_ _3349_/A _3349_/B vssd1 vssd1 vccd1 vccd1 _3351_/A sky130_fd_sc_hd__nand2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5019_ _5019_/CLK _5019_/D vssd1 vssd1 vccd1 vccd1 _5019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5189__96 vssd1 vssd1 vccd1 vccd1 _5189__96/HI _5297_/A sky130_fd_sc_hd__conb_1
XFILLER_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2720_ _2720_/A vssd1 vssd1 vccd1 vccd1 _4781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2651_ _4970_/Q _4762_/Q _2657_/S vssd1 vssd1 vccd1 vccd1 _2652_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2582_ _2592_/A _2582_/B vssd1 vssd1 vccd1 vccd1 _2583_/A sky130_fd_sc_hd__and2_1
X_4321_ _4321_/A vssd1 vssd1 vccd1 vccd1 _4321_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4252_ _4252_/A _4252_/B vssd1 vssd1 vccd1 vccd1 _4284_/A sky130_fd_sc_hd__nor2_1
X_3203_ _3203_/A _3203_/B vssd1 vssd1 vccd1 vccd1 _3233_/A sky130_fd_sc_hd__nor2_1
X_4183_ _5011_/Q _4791_/Q vssd1 vssd1 vccd1 vccd1 _4189_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3134_ _4022_/A vssd1 vssd1 vccd1 vccd1 _3551_/A sky130_fd_sc_hd__clkbuf_2
X_3065_ _3046_/A _3048_/Y _3053_/B _3061_/A _3051_/Y vssd1 vssd1 vccd1 vccd1 _3065_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3967_ _4983_/Q _4763_/Q vssd1 vssd1 vccd1 vccd1 _3967_/X sky130_fd_sc_hd__or2_1
XFILLER_10_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2918_ _2918_/A vssd1 vssd1 vccd1 vccd1 _4832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3898_ _3895_/Y _3889_/X _3901_/B _3903_/C vssd1 vssd1 vccd1 vccd1 _3898_/Y sky130_fd_sc_hd__a22oi_1
X_2849_ _2849_/A vssd1 vssd1 vccd1 vccd1 _4818_/D sky130_fd_sc_hd__clkbuf_1
X_4519_ _4522_/A _4519_/B vssd1 vssd1 vccd1 vccd1 _4520_/A sky130_fd_sc_hd__and2_1
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4870_ _5050_/CLK _4870_/D vssd1 vssd1 vccd1 vccd1 _4870_/Q sky130_fd_sc_hd__dfxtp_1
X_3821_ _3819_/Y _3821_/B vssd1 vssd1 vccd1 vccd1 _3821_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3752_ _4957_/Q _4737_/Q vssd1 vssd1 vccd1 vccd1 _3754_/B sky130_fd_sc_hd__xnor2_1
X_2703_ _4985_/Q _4777_/Q _2710_/S vssd1 vssd1 vccd1 vccd1 _2704_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3683_ _5116_/Q _4948_/Q vssd1 vssd1 vccd1 vccd1 _3685_/A sky130_fd_sc_hd__and2_1
X_2634_ _2645_/A _2634_/B vssd1 vssd1 vccd1 vccd1 _2635_/A sky130_fd_sc_hd__and2_1
X_2565_ _2575_/A _2565_/B vssd1 vssd1 vccd1 vccd1 _2566_/A sky130_fd_sc_hd__and2_1
X_4304_ _4290_/A _4292_/Y _4297_/B _4295_/Y vssd1 vssd1 vccd1 vccd1 _4305_/B sky130_fd_sc_hd__a31o_1
X_2496_ _2497_/A vssd1 vssd1 vccd1 vccd1 _2496_/Y sky130_fd_sc_hd__inv_2
X_5284_ _5284_/A _2480_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
X_4235_ _5017_/Q _4797_/Q vssd1 vssd1 vccd1 vccd1 _4235_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4166_ _4190_/A _4161_/B _4157_/A vssd1 vssd1 vccd1 vccd1 _4170_/A sky130_fd_sc_hd__a21oi_1
XFILLER_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3117_ _3116_/A _3138_/B _3084_/X vssd1 vssd1 vccd1 vccd1 _3117_/X sky130_fd_sc_hd__a21o_1
X_4097_ _4999_/Q _4779_/Q _4095_/Y _4093_/C _4096_/X vssd1 vssd1 vccd1 vccd1 _4097_/X
+ sky130_fd_sc_hd__a221o_1
X_3048_ _3048_/A _3048_/B vssd1 vssd1 vccd1 vccd1 _3048_/Y sky130_fd_sc_hd__nand2_1
X_4999_ _4999_/CLK _4999_/D vssd1 vssd1 vccd1 vccd1 _4999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5159__66 vssd1 vssd1 vccd1 vccd1 _5159__66/HI _5254_/A sky130_fd_sc_hd__conb_1
XFILLER_9_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4975_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5173__80 vssd1 vssd1 vccd1 vccd1 _5173__80/HI _5268_/A sky130_fd_sc_hd__conb_1
X_4020_ _4020_/A _4020_/B vssd1 vssd1 vccd1 vccd1 _4020_/Y sky130_fd_sc_hd__xnor2_1
X_4922_ _5103_/CLK _4922_/D vssd1 vssd1 vccd1 vccd1 _4922_/Q sky130_fd_sc_hd__dfxtp_1
X_4853_ _5032_/CLK _4853_/D vssd1 vssd1 vccd1 vccd1 _4853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4784_ _5004_/CLK _4784_/D vssd1 vssd1 vccd1 vccd1 _4784_/Q sky130_fd_sc_hd__dfxtp_1
X_3804_ _4951_/Q _3784_/X _3802_/Y _3803_/X _3773_/X vssd1 vssd1 vccd1 vccd1 _4951_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3735_ _3720_/A _3722_/Y _3728_/B _3726_/Y vssd1 vssd1 vccd1 vccd1 _3736_/B sky130_fd_sc_hd__a31o_1
X_3666_ _4934_/Q vssd1 vssd1 vccd1 vccd1 _3666_/Y sky130_fd_sc_hd__inv_2
X_2617_ _2627_/A _2617_/B vssd1 vssd1 vccd1 vccd1 _2618_/A sky130_fd_sc_hd__and2_1
X_3597_ _3597_/A _3597_/B vssd1 vssd1 vccd1 vccd1 _3617_/B sky130_fd_sc_hd__and2_1
X_2548_ _2548_/A vssd1 vssd1 vccd1 vccd1 _2548_/Y sky130_fd_sc_hd__inv_2
X_5267_ _5267_/A _2458_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
X_4218_ _5003_/Q _4165_/X _4216_/X _4217_/Y _4187_/X vssd1 vssd1 vccd1 vccd1 _5003_/D
+ sky130_fd_sc_hd__o221a_1
X_2479_ _2485_/A vssd1 vssd1 vccd1 vccd1 _2484_/A sky130_fd_sc_hd__clkbuf_16
X_4149_ _5007_/Q _4787_/Q vssd1 vssd1 vccd1 vccd1 _4151_/A sky130_fd_sc_hd__nor2_1
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3520_ _3520_/A _3521_/C vssd1 vssd1 vccd1 vccd1 _3529_/A sky130_fd_sc_hd__or2_1
X_3451_ _4919_/Q _5087_/Q vssd1 vssd1 vccd1 vccd1 _3451_/Y sky130_fd_sc_hd__xnor2_1
X_3382_ _3383_/A _3383_/B vssd1 vssd1 vccd1 vccd1 _3382_/X sky130_fd_sc_hd__or2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5121_ _5121_/CLK _5121_/D vssd1 vssd1 vccd1 vccd1 _5121_/Q sky130_fd_sc_hd__dfxtp_1
X_5052_ _5058_/CLK _5052_/D vssd1 vssd1 vccd1 vccd1 _5052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4003_ _4003_/A _4003_/B vssd1 vssd1 vccd1 vccd1 _4004_/C sky130_fd_sc_hd__nand2_1
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4905_ _5094_/CLK _4905_/D vssd1 vssd1 vccd1 vccd1 _4905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4836_ _4836_/CLK _4836_/D vssd1 vssd1 vccd1 vccd1 _5277_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4767_ _4975_/CLK _4767_/D vssd1 vssd1 vccd1 vccd1 _4767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5129__36 vssd1 vssd1 vccd1 vccd1 _5129__36/HI _5224_/A sky130_fd_sc_hd__conb_1
X_4698_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__clkbuf_2
X_3718_ _5120_/Q _4952_/Q vssd1 vssd1 vccd1 vccd1 _3720_/A sky130_fd_sc_hd__nand2_1
X_3649_ _3936_/B vssd1 vssd1 vccd1 vccd1 _3931_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5319_ _5319_/A _2521_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
XFILLER_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5143__50 vssd1 vssd1 vccd1 vccd1 _5143__50/HI _5238_/A sky130_fd_sc_hd__conb_1
XFILLER_10_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2951_ _2951_/A _2951_/B vssd1 vssd1 vccd1 vccd1 _2952_/A sky130_fd_sc_hd__and2_1
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5094_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4621_ _4621_/A vssd1 vssd1 vccd1 vccd1 _5089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2882_ _2862_/X input8/X _2863_/X vssd1 vssd1 vccd1 vccd1 _2882_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4552_ _4552_/A vssd1 vssd1 vccd1 vccd1 _5069_/D sky130_fd_sc_hd__clkbuf_1
X_3503_ _3566_/A vssd1 vssd1 vccd1 vccd1 _3503_/X sky130_fd_sc_hd__clkbuf_2
X_4483_ _4483_/A vssd1 vssd1 vccd1 vccd1 _5049_/D sky130_fd_sc_hd__clkbuf_1
X_3434_ _3566_/A vssd1 vssd1 vccd1 vccd1 _3434_/X sky130_fd_sc_hd__clkbuf_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _4908_/Q _5076_/Q vssd1 vssd1 vccd1 vccd1 _3372_/A sky130_fd_sc_hd__nand2_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _4887_/Q _3268_/X _3294_/Y _3295_/X _3230_/X vssd1 vssd1 vccd1 vccd1 _4887_/D
+ sky130_fd_sc_hd__o221a_1
X_5104_ _5106_/CLK _5104_/D vssd1 vssd1 vccd1 vccd1 _5104_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5046_/CLK _5035_/D vssd1 vssd1 vccd1 vccd1 _5035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4819_ _5027_/CLK _4819_/D vssd1 vssd1 vccd1 vccd1 _4819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3150_ _4881_/Q _5049_/Q vssd1 vssd1 vccd1 vccd1 _3150_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3081_ _4873_/Q _5041_/Q vssd1 vssd1 vccd1 vccd1 _3083_/B sky130_fd_sc_hd__xnor2_1
X_3983_ _3996_/A _3984_/B vssd1 vssd1 vccd1 vccd1 _3983_/X sky130_fd_sc_hd__or2_1
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2934_ _2934_/A _2934_/B vssd1 vssd1 vccd1 vccd1 _2935_/A sky130_fd_sc_hd__and2_1
X_2865_ _2889_/A vssd1 vssd1 vccd1 vccd1 _2865_/X sky130_fd_sc_hd__clkbuf_2
X_4604_ _4604_/A vssd1 vssd1 vccd1 vccd1 _5084_/D sky130_fd_sc_hd__clkbuf_1
X_4535_ _4885_/Q _5065_/Q _4542_/S vssd1 vssd1 vccd1 vccd1 _4536_/B sky130_fd_sc_hd__mux2_1
X_2796_ _2803_/A _2796_/B vssd1 vssd1 vccd1 vccd1 _2797_/A sky130_fd_sc_hd__and2_1
X_4466_ _4865_/Q _5045_/Q _4474_/S vssd1 vssd1 vccd1 vccd1 _4467_/B sky130_fd_sc_hd__mux2_1
X_3417_ _4914_/Q _5082_/Q _3421_/A _3412_/B vssd1 vssd1 vccd1 vccd1 _3417_/Y sky130_fd_sc_hd__a22oi_1
X_4397_ _4397_/A _4397_/B vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__or2_1
X_3348_ _4906_/Q _5074_/Q vssd1 vssd1 vccd1 vccd1 _3349_/B sky130_fd_sc_hd__nand2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _3566_/A vssd1 vssd1 vccd1 vccd1 _3279_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5018_ _5018_/CLK _5018_/D vssd1 vssd1 vccd1 vccd1 _5018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2650_ _2650_/A vssd1 vssd1 vccd1 vccd1 _4761_/D sky130_fd_sc_hd__clkbuf_1
X_2581_ _4950_/Q _4742_/Q _2587_/S vssd1 vssd1 vccd1 vccd1 _2582_/B sky130_fd_sc_hd__mux2_1
X_4320_ _4316_/X _4325_/A _4319_/X vssd1 vssd1 vccd1 vccd1 _4320_/X sky130_fd_sc_hd__a21o_1
X_4251_ _5020_/Q _4800_/Q vssd1 vssd1 vccd1 vccd1 _4252_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3202_ _4888_/Q _5056_/Q vssd1 vssd1 vccd1 vccd1 _3203_/B sky130_fd_sc_hd__nor2_1
X_4182_ _5010_/Q _4790_/Q vssd1 vssd1 vccd1 vccd1 _4182_/Y sky130_fd_sc_hd__nand2_1
X_3133_ _3133_/A vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__clkbuf_2
X_3064_ _2980_/X _3061_/X _3062_/X _3063_/X vssd1 vssd1 vccd1 vccd1 _4858_/D sky130_fd_sc_hd__o211a_1
X_3966_ _3966_/A _3966_/B vssd1 vssd1 vccd1 vccd1 _3971_/A sky130_fd_sc_hd__nor2_1
X_2917_ _2917_/A _2917_/B vssd1 vssd1 vccd1 vccd1 _2918_/A sky130_fd_sc_hd__and2_1
X_3897_ _4975_/Q _4755_/Q vssd1 vssd1 vccd1 vccd1 _3903_/C sky130_fd_sc_hd__or2_1
X_2848_ _2917_/A _2848_/B vssd1 vssd1 vccd1 vccd1 _2849_/A sky130_fd_sc_hd__and2_1
X_2779_ _5007_/Q _4799_/Q _2779_/S vssd1 vssd1 vccd1 vccd1 _2780_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4518_ _4880_/Q _5060_/Q _4525_/S vssd1 vssd1 vccd1 vccd1 _4519_/B sky130_fd_sc_hd__mux2_1
X_4449_ _4452_/A _4449_/B vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__and2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3820_ _4965_/Q _4745_/Q vssd1 vssd1 vccd1 vccd1 _3821_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3751_ _4944_/Q _3745_/X _3750_/X _3724_/X vssd1 vssd1 vccd1 vccd1 _4944_/D sky130_fd_sc_hd__o211a_1
X_2702_ _2702_/A vssd1 vssd1 vccd1 vccd1 _4776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3682_ _4935_/Q _3664_/A _3679_/Y _3681_/X _3646_/X vssd1 vssd1 vccd1 vccd1 _4935_/D
+ sky130_fd_sc_hd__o221a_1
X_2633_ _4965_/Q _4757_/Q _2639_/S vssd1 vssd1 vccd1 vccd1 _2634_/B sky130_fd_sc_hd__mux2_1
X_2564_ _4945_/Q _4737_/Q _2570_/S vssd1 vssd1 vccd1 vccd1 _2565_/B sky130_fd_sc_hd__mux2_1
X_4303_ _4303_/A _4303_/B vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__or2_1
X_5283_ _5283_/A _2478_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
X_2495_ _2497_/A vssd1 vssd1 vccd1 vccd1 _2495_/Y sky130_fd_sc_hd__inv_2
X_4234_ _5006_/Q vssd1 vssd1 vccd1 vccd1 _4234_/Y sky130_fd_sc_hd__inv_2
X_4165_ _4212_/B vssd1 vssd1 vccd1 vccd1 _4165_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3116_ _3116_/A _3138_/B vssd1 vssd1 vccd1 vccd1 _3116_/Y sky130_fd_sc_hd__nor2_1
X_4096_ _4998_/Q _4778_/Q _4096_/C vssd1 vssd1 vccd1 vccd1 _4096_/X sky130_fd_sc_hd__and3_1
XFILLER_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3047_ _3048_/A _3048_/B vssd1 vssd1 vccd1 vccd1 _3047_/X sky130_fd_sc_hd__or2_1
XFILLER_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4998_ _5002_/CLK _4998_/D vssd1 vssd1 vccd1 vccd1 _4998_/Q sky130_fd_sc_hd__dfxtp_2
X_3949_ _3942_/A _3942_/B _3948_/Y vssd1 vssd1 vccd1 vccd1 _3954_/A sky130_fd_sc_hd__o21ai_1
XFILLER_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4921_ _5103_/CLK _4921_/D vssd1 vssd1 vccd1 vccd1 _4921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4852_ _5041_/CLK _4852_/D vssd1 vssd1 vccd1 vccd1 _4852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3803_ _3805_/B _3805_/C _3801_/Y _3755_/A vssd1 vssd1 vccd1 vccd1 _3803_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4783_ _5004_/CLK _4783_/D vssd1 vssd1 vccd1 vccd1 _4783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3734_ _3734_/A _3734_/B vssd1 vssd1 vccd1 vccd1 _3736_/A sky130_fd_sc_hd__or2_1
X_3665_ _4933_/Q _3652_/X _3664_/Y _3659_/X vssd1 vssd1 vccd1 vccd1 _4933_/D sky130_fd_sc_hd__o211a_1
X_2616_ _4960_/Q _4752_/Q _2622_/S vssd1 vssd1 vccd1 vccd1 _2617_/B sky130_fd_sc_hd__mux2_1
X_3596_ _4937_/Q _5105_/Q vssd1 vssd1 vccd1 vccd1 _3597_/B sky130_fd_sc_hd__nand2_1
X_2547_ _2548_/A vssd1 vssd1 vccd1 vccd1 _2547_/Y sky130_fd_sc_hd__inv_2
X_2478_ _2478_/A vssd1 vssd1 vccd1 vccd1 _2478_/Y sky130_fd_sc_hd__inv_2
X_5266_ _5266_/A _2457_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
X_4217_ _4209_/B _4214_/Y _4215_/Y _4165_/X vssd1 vssd1 vccd1 vccd1 _4217_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4148_ _4139_/Y _4130_/X _4147_/Y _3360_/X vssd1 vssd1 vccd1 vccd1 _4994_/D sky130_fd_sc_hd__a211oi_1
XFILLER_83_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _4074_/A _4073_/B _4071_/Y vssd1 vssd1 vccd1 vccd1 _4086_/B sky130_fd_sc_hd__a21o_1
X_5194__101 vssd1 vssd1 vccd1 vccd1 _5194__101/HI _5302_/A sky130_fd_sc_hd__conb_1
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3450_ _3430_/A _3432_/Y _3438_/B _3447_/A _3436_/Y vssd1 vssd1 vccd1 vccd1 _3450_/Y
+ sky130_fd_sc_hd__a311oi_2
X_3381_ _3381_/A _3381_/B vssd1 vssd1 vccd1 vccd1 _3383_/B sky130_fd_sc_hd__and2_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5120_ _5121_/CLK _5120_/D vssd1 vssd1 vccd1 vccd1 _5120_/Q sky130_fd_sc_hd__dfxtp_1
X_5051_ _5051_/CLK _5051_/D vssd1 vssd1 vccd1 vccd1 _5051_/Q sky130_fd_sc_hd__dfxtp_1
X_4002_ _4988_/Q _4768_/Q vssd1 vssd1 vccd1 vccd1 _4003_/B sky130_fd_sc_hd__or2_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4904_ _5085_/CLK _4904_/D vssd1 vssd1 vccd1 vccd1 _4904_/Q sky130_fd_sc_hd__dfxtp_1
X_4835_ _5033_/CLK _4835_/D vssd1 vssd1 vccd1 vccd1 _5276_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4766_ _4989_/CLK _4766_/D vssd1 vssd1 vccd1 vccd1 _4766_/Q sky130_fd_sc_hd__dfxtp_1
X_3717_ _3689_/B _3712_/X _3716_/X vssd1 vssd1 vccd1 vccd1 _3722_/A sky130_fd_sc_hd__a21o_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4697_ _4697_/A vssd1 vssd1 vccd1 vccd1 _5111_/D sky130_fd_sc_hd__clkbuf_1
X_3648_ _3648_/A _4030_/B vssd1 vssd1 vccd1 vccd1 _3936_/B sky130_fd_sc_hd__or2b_1
X_3579_ _4935_/Q _5103_/Q vssd1 vssd1 vccd1 vccd1 _3580_/B sky130_fd_sc_hd__and2_1
X_5318_ _5318_/A _2520_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
X_5249_ _5249_/A _2548_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
Xclkbuf_leaf_2_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5050_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2950_ _5283_/A _4858_/Q _2954_/S vssd1 vssd1 vccd1 vccd1 _2951_/B sky130_fd_sc_hd__mux2_1
X_2881_ _2878_/X _4824_/Q _2879_/X _2880_/X _2876_/X vssd1 vssd1 vccd1 vccd1 _4824_/D
+ sky130_fd_sc_hd__o221a_1
X_4620_ _4626_/A _4620_/B vssd1 vssd1 vccd1 vccd1 _4621_/A sky130_fd_sc_hd__and2_1
XFILLER_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4551_ _4557_/A _4551_/B vssd1 vssd1 vccd1 vccd1 _4552_/A sky130_fd_sc_hd__and2_1
X_3502_ _4913_/Q _3544_/B vssd1 vssd1 vccd1 vccd1 _3502_/X sky130_fd_sc_hd__or2_1
X_4482_ _4488_/A _4482_/B vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__and2_1
X_3433_ _3431_/X _3432_/Y _3373_/X vssd1 vssd1 vccd1 vccd1 _3433_/X sky130_fd_sc_hd__a21o_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _4908_/Q _5076_/Q vssd1 vssd1 vccd1 vccd1 _3364_/X sky130_fd_sc_hd__or2_1
X_5103_ _5103_/CLK _5103_/D vssd1 vssd1 vccd1 vccd1 _5103_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3285_/A _3287_/Y _3293_/Y _3288_/X vssd1 vssd1 vccd1 vccd1 _3295_/X sky130_fd_sc_hd__a31o_1
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5046_/CLK _5034_/D vssd1 vssd1 vccd1 vccd1 _5034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4818_ _5027_/CLK _4818_/D vssd1 vssd1 vccd1 vccd1 _4818_/Q sky130_fd_sc_hd__dfxtp_1
X_4749_ _4752_/CLK _4749_/D vssd1 vssd1 vccd1 vccd1 _4749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3080_ _4860_/Q _3074_/X _3079_/X _3063_/X vssd1 vssd1 vccd1 vccd1 _4860_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3982_ _3978_/A _3976_/Y _3977_/A vssd1 vssd1 vccd1 vccd1 _3984_/B sky130_fd_sc_hd__a21o_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2933_ _5278_/A _4853_/Q _2944_/S vssd1 vssd1 vccd1 vccd1 _2934_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2864_ _2862_/X input4/X _2863_/X vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__o21a_1
X_4603_ _4609_/A _4603_/B vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__and2_1
X_2795_ _5011_/Q _4803_/Q _2798_/S vssd1 vssd1 vccd1 vccd1 _2796_/B sky130_fd_sc_hd__mux2_1
X_4534_ _4534_/A vssd1 vssd1 vccd1 vccd1 _5064_/D sky130_fd_sc_hd__clkbuf_1
X_4465_ _4465_/A vssd1 vssd1 vccd1 vccd1 _5044_/D sky130_fd_sc_hd__clkbuf_1
X_3416_ _4915_/Q _5083_/Q vssd1 vssd1 vccd1 vccd1 _3421_/C sky130_fd_sc_hd__or2_1
X_4396_ _4830_/Q _4818_/Q vssd1 vssd1 vccd1 vccd1 _4397_/B sky130_fd_sc_hd__and2_1
X_3347_ _4906_/Q _5074_/Q vssd1 vssd1 vccd1 vccd1 _3349_/A sky130_fd_sc_hd__or2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _4022_/A vssd1 vssd1 vccd1 vccd1 _3566_/A sky130_fd_sc_hd__buf_2
X_5017_ _5018_/CLK _5017_/D vssd1 vssd1 vccd1 vccd1 _5017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2580_ _2580_/A vssd1 vssd1 vccd1 vccd1 _4741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _5020_/Q _4800_/Q vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__and2_1
XFILLER_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4181_ _4998_/Q _4126_/X _4180_/X _4163_/X vssd1 vssd1 vccd1 vccd1 _4998_/D sky130_fd_sc_hd__o211a_1
X_3201_ _4888_/Q _5056_/Q vssd1 vssd1 vccd1 vccd1 _3203_/A sky130_fd_sc_hd__and2_1
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3132_ _3128_/Y _3122_/X _3137_/B _3139_/C _3084_/A vssd1 vssd1 vccd1 vccd1 _3132_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_82_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3063_ _4733_/A vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3965_ _4984_/Q _4764_/Q vssd1 vssd1 vccd1 vccd1 _3966_/B sky130_fd_sc_hd__nor2_1
X_3896_ _4975_/Q _4755_/Q vssd1 vssd1 vccd1 vccd1 _3901_/B sky130_fd_sc_hd__nand2_1
X_2916_ _5273_/A _4848_/Q _2968_/B vssd1 vssd1 vccd1 vccd1 _2917_/B sky130_fd_sc_hd__mux2_1
X_2847_ _5026_/Q _4818_/Q _2850_/S vssd1 vssd1 vccd1 vccd1 _2848_/B sky130_fd_sc_hd__mux2_1
X_2778_ _2778_/A vssd1 vssd1 vccd1 vccd1 _4798_/D sky130_fd_sc_hd__clkbuf_1
X_4517_ _4517_/A vssd1 vssd1 vccd1 vccd1 _5059_/D sky130_fd_sc_hd__clkbuf_1
X_4448_ _4860_/Q _5040_/Q _4455_/S vssd1 vssd1 vccd1 vccd1 _4449_/B sky130_fd_sc_hd__mux2_1
X_4379_ _4826_/Q _4814_/Q _4379_/C vssd1 vssd1 vccd1 vccd1 _4379_/X sky130_fd_sc_hd__and3_1
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3750_ _3746_/X _3754_/A _3749_/X vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__a21o_1
X_2701_ _2715_/A _2701_/B vssd1 vssd1 vccd1 vccd1 _2702_/A sky130_fd_sc_hd__and2_1
XFILLER_9_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3681_ _3671_/A _3673_/Y _3678_/Y _3680_/X vssd1 vssd1 vccd1 vccd1 _3681_/X sky130_fd_sc_hd__a31o_1
X_2632_ _2632_/A vssd1 vssd1 vccd1 vccd1 _4756_/D sky130_fd_sc_hd__clkbuf_1
X_2563_ _2563_/A vssd1 vssd1 vccd1 vccd1 _4736_/D sky130_fd_sc_hd__clkbuf_1
X_5282_ _5282_/A _2477_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
X_4302_ _5026_/Q _4806_/Q vssd1 vssd1 vccd1 vccd1 _4303_/B sky130_fd_sc_hd__and2_1
X_2494_ _2497_/A vssd1 vssd1 vccd1 vccd1 _2494_/Y sky130_fd_sc_hd__inv_2
X_4233_ _5005_/Q _4220_/X _4231_/X _4232_/X vssd1 vssd1 vccd1 vccd1 _5005_/D sky130_fd_sc_hd__o211a_1
X_4164_ _4130_/X _4161_/X _4162_/X _4163_/X vssd1 vssd1 vccd1 vccd1 _4996_/D sky130_fd_sc_hd__o211a_1
X_4095_ _4094_/Y _4073_/B _4071_/Y vssd1 vssd1 vccd1 vccd1 _4095_/Y sky130_fd_sc_hd__a21oi_1
X_3115_ _3115_/A _3115_/B vssd1 vssd1 vccd1 vccd1 _3138_/B sky130_fd_sc_hd__and2_1
XFILLER_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3046_ _3046_/A _3046_/B vssd1 vssd1 vccd1 vccd1 _3048_/B sky130_fd_sc_hd__and2_1
X_4997_ _5002_/CLK _4997_/D vssd1 vssd1 vccd1 vccd1 _4997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3948_ _4981_/Q _4761_/Q vssd1 vssd1 vccd1 vccd1 _3948_/Y sky130_fd_sc_hd__nand2_1
X_3879_ _3902_/A _3874_/B _3870_/A vssd1 vssd1 vccd1 vccd1 _3883_/A sky130_fd_sc_hd__a21oi_1
XFILLER_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4954_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4920_ _5101_/CLK _4920_/D vssd1 vssd1 vccd1 vccd1 _4920_/Q sky130_fd_sc_hd__dfxtp_1
X_4851_ _5033_/CLK _4851_/D vssd1 vssd1 vccd1 vccd1 _4851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3802_ _3805_/B _3805_/C _3801_/Y vssd1 vssd1 vccd1 vccd1 _3802_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4782_ _5004_/CLK _4782_/D vssd1 vssd1 vccd1 vccd1 _4782_/Q sky130_fd_sc_hd__dfxtp_1
X_3733_ _5122_/Q _4954_/Q vssd1 vssd1 vccd1 vccd1 _3734_/B sky130_fd_sc_hd__and2_1
X_3664_ _3664_/A _3664_/B vssd1 vssd1 vccd1 vccd1 _3664_/Y sky130_fd_sc_hd__nand2_1
X_2615_ _2615_/A vssd1 vssd1 vccd1 vccd1 _4751_/D sky130_fd_sc_hd__clkbuf_1
X_3595_ _4937_/Q _5105_/Q vssd1 vssd1 vccd1 vccd1 _3597_/A sky130_fd_sc_hd__or2_1
X_2546_ _2548_/A vssd1 vssd1 vccd1 vccd1 _2546_/Y sky130_fd_sc_hd__inv_2
X_5164__71 vssd1 vssd1 vccd1 vccd1 _5164__71/HI _5259_/A sky130_fd_sc_hd__conb_1
X_5265_ _5265_/A _2456_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
X_2477_ _2478_/A vssd1 vssd1 vccd1 vccd1 _2477_/Y sky130_fd_sc_hd__inv_2
X_4216_ _4209_/B _4214_/Y _4215_/Y vssd1 vssd1 vccd1 vccd1 _4216_/X sky130_fd_sc_hd__o21a_1
X_4147_ _4145_/X _4146_/Y _4130_/X vssd1 vssd1 vccd1 vccd1 _4147_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4078_ _4998_/Q _4778_/Q vssd1 vssd1 vccd1 vccd1 _4092_/A sky130_fd_sc_hd__xor2_2
XFILLER_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3029_ _3040_/A _3013_/B _3019_/A _3039_/A _3028_/Y vssd1 vssd1 vccd1 vccd1 _3029_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3380_ _4910_/Q _5078_/Q vssd1 vssd1 vccd1 vccd1 _3381_/B sky130_fd_sc_hd__or2_1
XFILLER_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _5050_/CLK _5050_/D vssd1 vssd1 vccd1 vccd1 _5050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4001_ _4988_/Q _4768_/Q vssd1 vssd1 vccd1 vccd1 _4003_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4903_ _5085_/CLK _4903_/D vssd1 vssd1 vccd1 vccd1 _4903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4834_ _4836_/CLK _4834_/D vssd1 vssd1 vccd1 vccd1 _5275_/A sky130_fd_sc_hd__dfxtp_1
X_4765_ _4981_/CLK _4765_/D vssd1 vssd1 vccd1 vccd1 _4765_/Q sky130_fd_sc_hd__dfxtp_1
X_3716_ _3714_/Y _3712_/C _3715_/X _3711_/C vssd1 vssd1 vccd1 vccd1 _3716_/X sky130_fd_sc_hd__a22o_1
X_4696_ _4696_/A _4696_/B vssd1 vssd1 vccd1 vccd1 _4697_/A sky130_fd_sc_hd__and2_1
X_3647_ _4931_/Q _3593_/X _3643_/X _3644_/Y _3646_/X vssd1 vssd1 vccd1 vccd1 _4931_/D
+ sky130_fd_sc_hd__o221a_1
X_3578_ _4935_/Q _5103_/Q vssd1 vssd1 vccd1 vccd1 _3580_/A sky130_fd_sc_hd__nor2_1
X_2529_ _2533_/A vssd1 vssd1 vccd1 vccd1 _2529_/Y sky130_fd_sc_hd__inv_2
X_5317_ _5317_/A _2519_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
X_5248_ _5248_/A _2547_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2880_ _2865_/X input22/X _2878_/A vssd1 vssd1 vccd1 vccd1 _2880_/X sky130_fd_sc_hd__a21bo_1
X_4550_ _4889_/Q _5069_/Q _4561_/S vssd1 vssd1 vccd1 vccd1 _4551_/B sky130_fd_sc_hd__mux2_1
X_3501_ _3501_/A _3522_/A vssd1 vssd1 vccd1 vccd1 _3501_/X sky130_fd_sc_hd__xor2_1
X_4481_ _4869_/Q _5049_/Q _4491_/S vssd1 vssd1 vccd1 vccd1 _4482_/B sky130_fd_sc_hd__mux2_1
X_3432_ _3432_/A _3432_/B vssd1 vssd1 vccd1 vccd1 _3432_/Y sky130_fd_sc_hd__nand2_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _3448_/B vssd1 vssd1 vccd1 vccd1 _3363_/X sky130_fd_sc_hd__clkbuf_2
X_5134__41 vssd1 vssd1 vccd1 vccd1 _5134__41/HI _5229_/A sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5051_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5103_/CLK _5102_/D vssd1 vssd1 vccd1 vccd1 _5102_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _3285_/A _3287_/Y _3293_/Y vssd1 vssd1 vccd1 vccd1 _3294_/Y sky130_fd_sc_hd__a21oi_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/CLK _5033_/D vssd1 vssd1 vccd1 vccd1 _5033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4817_ _5027_/CLK _4817_/D vssd1 vssd1 vccd1 vccd1 _4817_/Q sky130_fd_sc_hd__dfxtp_1
X_4748_ _4964_/CLK _4748_/D vssd1 vssd1 vccd1 vccd1 _4748_/Q sky130_fd_sc_hd__dfxtp_1
X_4679_ _4679_/A _4679_/B vssd1 vssd1 vccd1 vccd1 _4680_/A sky130_fd_sc_hd__and2_1
XFILLER_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3981_ _4986_/Q _4766_/Q vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__xnor2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2932_ _2932_/A vssd1 vssd1 vccd1 vccd1 _4836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2863_ _2905_/A vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4602_ _4904_/Q _5084_/Q _4612_/S vssd1 vssd1 vccd1 vccd1 _4603_/B sky130_fd_sc_hd__mux2_1
X_2794_ _2794_/A vssd1 vssd1 vccd1 vccd1 _4802_/D sky130_fd_sc_hd__clkbuf_1
X_4533_ _4539_/A _4533_/B vssd1 vssd1 vccd1 vccd1 _4534_/A sky130_fd_sc_hd__and2_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ _4470_/A _4464_/B vssd1 vssd1 vccd1 vccd1 _4465_/A sky130_fd_sc_hd__and2_1
X_3415_ _4915_/Q _5083_/Q vssd1 vssd1 vccd1 vccd1 _3421_/B sky130_fd_sc_hd__nand2_1
X_4395_ _4830_/Q _4818_/Q vssd1 vssd1 vccd1 vccd1 _4397_/A sky130_fd_sc_hd__nor2_1
X_3346_ _4893_/Q _3277_/A _3344_/Y _3345_/X _3325_/X vssd1 vssd1 vccd1 vccd1 _4893_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3277_/A _3277_/B vssd1 vssd1 vccd1 vccd1 _3277_/Y sky130_fd_sc_hd__nand2_1
X_5016_ _5018_/CLK _5016_/D vssd1 vssd1 vccd1 vccd1 _5016_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4180_ _4176_/X _4179_/X _4136_/X vssd1 vssd1 vccd1 vccd1 _4180_/X sky130_fd_sc_hd__a21o_1
X_3200_ _4875_/Q _3172_/X _3198_/Y _3199_/X _3135_/X vssd1 vssd1 vccd1 vccd1 _4875_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3131_ _3128_/Y _3122_/X _3137_/B _3139_/C vssd1 vssd1 vccd1 vccd1 _3131_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3062_ _4858_/Q _3062_/B vssd1 vssd1 vccd1 vccd1 _3062_/X sky130_fd_sc_hd__or2_1
XFILLER_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ _4984_/Q _4764_/Q vssd1 vssd1 vccd1 vccd1 _3966_/A sky130_fd_sc_hd__and2_1
X_3895_ _4974_/Q _4754_/Q vssd1 vssd1 vccd1 vccd1 _3895_/Y sky130_fd_sc_hd__nand2_1
X_2915_ _2954_/S vssd1 vssd1 vccd1 vccd1 _2968_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2846_ _2846_/A vssd1 vssd1 vccd1 vccd1 _4817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2777_ _2784_/A _2777_/B vssd1 vssd1 vccd1 vccd1 _2778_/A sky130_fd_sc_hd__and2_1
X_4516_ _4522_/A _4516_/B vssd1 vssd1 vccd1 vccd1 _4517_/A sky130_fd_sc_hd__and2_1
X_4447_ _4447_/A vssd1 vssd1 vccd1 vccd1 _5039_/D sky130_fd_sc_hd__clkbuf_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4378_ _4377_/Y _4357_/B _4355_/Y vssd1 vssd1 vccd1 vccd1 _4378_/Y sky130_fd_sc_hd__a21oi_1
X_3329_ _4900_/Q _5068_/Q vssd1 vssd1 vccd1 vccd1 _3329_/Y sky130_fd_sc_hd__nand2_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2700_ _4984_/Q _4776_/Q _2710_/S vssd1 vssd1 vccd1 vccd1 _2701_/B sky130_fd_sc_hd__mux2_1
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3680_ _3680_/A vssd1 vssd1 vccd1 vccd1 _3680_/X sky130_fd_sc_hd__clkbuf_2
X_2631_ _2645_/A _2631_/B vssd1 vssd1 vccd1 vccd1 _2632_/A sky130_fd_sc_hd__and2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2562_ _2575_/A _2562_/B vssd1 vssd1 vccd1 vccd1 _2563_/A sky130_fd_sc_hd__and2_1
X_5281_ _5281_/A _2476_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
X_4301_ _5026_/Q _4806_/Q vssd1 vssd1 vccd1 vccd1 _4303_/A sky130_fd_sc_hd__nor2_1
X_2493_ _2497_/A vssd1 vssd1 vccd1 vccd1 _2493_/Y sky130_fd_sc_hd__inv_2
X_4232_ _4321_/A vssd1 vssd1 vccd1 vccd1 _4232_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4163_ _4321_/A vssd1 vssd1 vccd1 vccd1 _4163_/X sky130_fd_sc_hd__clkbuf_2
X_4094_ _4996_/Q _4776_/Q vssd1 vssd1 vccd1 vccd1 _4094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3114_ _4877_/Q _5045_/Q vssd1 vssd1 vccd1 vccd1 _3115_/B sky130_fd_sc_hd__nand2_1
X_3045_ _4868_/Q _5036_/Q vssd1 vssd1 vccd1 vccd1 _3046_/B sky130_fd_sc_hd__or2_1
XFILLER_82_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4996_ _5002_/CLK _4996_/D vssd1 vssd1 vccd1 vccd1 _4996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3947_ _4970_/Q vssd1 vssd1 vccd1 vccd1 _3947_/Y sky130_fd_sc_hd__inv_2
X_3878_ _3924_/B vssd1 vssd1 vccd1 vccd1 _3878_/X sky130_fd_sc_hd__clkbuf_2
X_2829_ _2829_/A vssd1 vssd1 vccd1 vccd1 _4812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _5030_/CLK _4850_/D vssd1 vssd1 vccd1 vccd1 _4850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3801_ _4962_/Q _4742_/Q _3805_/A _3795_/B vssd1 vssd1 vccd1 vccd1 _3801_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4781_ _5004_/CLK _4781_/D vssd1 vssd1 vccd1 vccd1 _4781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3732_ _5122_/Q _4954_/Q vssd1 vssd1 vccd1 vccd1 _3734_/A sky130_fd_sc_hd__nor2_1
X_3663_ _3663_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3664_/B sky130_fd_sc_hd__xnor2_1
X_2614_ _2627_/A _2614_/B vssd1 vssd1 vccd1 vccd1 _2615_/A sky130_fd_sc_hd__and2_1
X_3594_ _3617_/A _3590_/B _3586_/A vssd1 vssd1 vccd1 vccd1 _3598_/A sky130_fd_sc_hd__a21oi_1
X_2545_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2545_/Y sky130_fd_sc_hd__inv_2
X_5264_ _5264_/A _2455_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
X_2476_ _2478_/A vssd1 vssd1 vccd1 vccd1 _2476_/Y sky130_fd_sc_hd__inv_2
X_4215_ _5015_/Q _4795_/Q vssd1 vssd1 vccd1 vccd1 _4215_/Y sky130_fd_sc_hd__xnor2_1
X_4146_ _4146_/A _4146_/B vssd1 vssd1 vccd1 vccd1 _4146_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4985_/Q _4043_/A _4074_/Y _4075_/X _4076_/X vssd1 vssd1 vccd1 vccd1 _4985_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3028_ _3027_/Y _3019_/B _3025_/Y vssd1 vssd1 vccd1 vccd1 _3028_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4979_ _5122_/CLK _4979_/D vssd1 vssd1 vccd1 vccd1 _4979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4000_ _3971_/A _3971_/B _3997_/Y _3999_/Y _3996_/B vssd1 vssd1 vccd1 vccd1 _4004_/B
+ sky130_fd_sc_hd__a311oi_2
XFILLER_1_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4902_ _5085_/CLK _4902_/D vssd1 vssd1 vccd1 vccd1 _4902_/Q sky130_fd_sc_hd__dfxtp_2
X_4833_ _5033_/CLK _4833_/D vssd1 vssd1 vccd1 vccd1 _5274_/A sky130_fd_sc_hd__dfxtp_1
X_4764_ _4966_/CLK _4764_/D vssd1 vssd1 vccd1 vccd1 _4764_/Q sky130_fd_sc_hd__dfxtp_1
X_3715_ _5119_/Q _4951_/Q _4950_/Q _5118_/Q vssd1 vssd1 vccd1 vccd1 _3715_/X sky130_fd_sc_hd__a22o_1
X_4695_ _4931_/Q _5111_/Q _4699_/S vssd1 vssd1 vccd1 vccd1 _4696_/B sky130_fd_sc_hd__mux2_1
X_3646_ _4076_/A vssd1 vssd1 vccd1 vccd1 _3646_/X sky130_fd_sc_hd__buf_2
X_3577_ _3568_/Y _3558_/X _3576_/Y _3479_/X vssd1 vssd1 vccd1 vccd1 _4922_/D sky130_fd_sc_hd__a211oi_1
X_2528_ _2540_/A vssd1 vssd1 vccd1 vccd1 _2533_/A sky130_fd_sc_hd__buf_12
X_5316_ _5316_/A _2518_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
X_5247_ _5247_/A _2546_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
X_2459_ _2459_/A vssd1 vssd1 vccd1 vccd1 _2459_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4129_ _4129_/A _4223_/B vssd1 vssd1 vccd1 vccd1 _4136_/A sky130_fd_sc_hd__or2_2
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3500_ _3500_/A _3499_/Y vssd1 vssd1 vccd1 vccd1 _3522_/A sky130_fd_sc_hd__or2b_1
X_4480_ _4480_/A vssd1 vssd1 vccd1 vccd1 _5048_/D sky130_fd_sc_hd__clkbuf_1
X_3431_ _3432_/A _3432_/B vssd1 vssd1 vccd1 vccd1 _3431_/X sky130_fd_sc_hd__or2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _4125_/A _3553_/B vssd1 vssd1 vccd1 vccd1 _3448_/B sky130_fd_sc_hd__nor2_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5101_/CLK _5101_/D vssd1 vssd1 vccd1 vccd1 _5101_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3293_/A _3293_/B vssd1 vssd1 vccd1 vccd1 _3293_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5032_/CLK _5032_/D vssd1 vssd1 vccd1 vccd1 _5032_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4995_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4816_ _5027_/CLK _4816_/D vssd1 vssd1 vccd1 vccd1 _4816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4747_ _5122_/CLK _4747_/D vssd1 vssd1 vccd1 vccd1 _4747_/Q sky130_fd_sc_hd__dfxtp_1
X_4678_ _4926_/Q _5106_/Q _4682_/S vssd1 vssd1 vccd1 vccd1 _4679_/B sky130_fd_sc_hd__mux2_1
X_3629_ _4941_/Q _5109_/Q vssd1 vssd1 vccd1 vccd1 _3630_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5209__116 vssd1 vssd1 vccd1 vccd1 _5209__116/HI _5317_/A sky130_fd_sc_hd__conb_1
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3980_ _3937_/X _3978_/X _3979_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _4973_/D sky130_fd_sc_hd__o211a_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _2934_/A _2931_/B vssd1 vssd1 vccd1 vccd1 _2932_/A sky130_fd_sc_hd__and2_1
XFILLER_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4601_ _4601_/A vssd1 vssd1 vccd1 vccd1 _5083_/D sky130_fd_sc_hd__clkbuf_1
X_2862_ _2889_/A vssd1 vssd1 vccd1 vccd1 _2862_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2793_ _2803_/A _2793_/B vssd1 vssd1 vccd1 vccd1 _2794_/A sky130_fd_sc_hd__and2_1
X_4532_ _4884_/Q _5064_/Q _4542_/S vssd1 vssd1 vccd1 vccd1 _4533_/B sky130_fd_sc_hd__mux2_1
X_4463_ _4864_/Q _5044_/Q _4474_/S vssd1 vssd1 vccd1 vccd1 _4464_/B sky130_fd_sc_hd__mux2_1
X_3414_ _4902_/Q _3363_/X _3413_/X _3353_/X vssd1 vssd1 vccd1 vccd1 _4902_/D sky130_fd_sc_hd__o211a_1
X_4394_ _5025_/Q _4367_/A _4392_/Y _4393_/X _2557_/A vssd1 vssd1 vccd1 vccd1 _5025_/D
+ sky130_fd_sc_hd__o221a_1
X_3345_ _3336_/A _3338_/Y _3343_/X _3288_/A vssd1 vssd1 vccd1 vccd1 _3345_/X sky130_fd_sc_hd__a31o_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _3276_/A _3276_/B vssd1 vssd1 vccd1 vccd1 _3277_/B sky130_fd_sc_hd__xnor2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5015_/CLK _5015_/D vssd1 vssd1 vccd1 vccd1 _5015_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3130_ _4879_/Q _5047_/Q vssd1 vssd1 vccd1 vccd1 _3139_/C sky130_fd_sc_hd__or2_1
X_3061_ _3061_/A _3061_/B vssd1 vssd1 vccd1 vccd1 _3061_/X sky130_fd_sc_hd__xor2_1
XFILLER_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3963_ _4971_/Q _3933_/A _3960_/Y _3961_/X _3962_/X vssd1 vssd1 vccd1 vccd1 _4971_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_16_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3894_ _4962_/Q _3838_/X _3893_/X _3876_/X vssd1 vssd1 vccd1 vccd1 _4962_/D sky130_fd_sc_hd__o211a_1
X_2914_ _3648_/A _2967_/B vssd1 vssd1 vccd1 vccd1 _2954_/S sky130_fd_sc_hd__and2_2
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2845_ _2917_/A _2845_/B vssd1 vssd1 vccd1 vccd1 _2846_/A sky130_fd_sc_hd__and2_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4515_ _4879_/Q _5059_/Q _4525_/S vssd1 vssd1 vccd1 vccd1 _4516_/B sky130_fd_sc_hd__mux2_1
X_2776_ _5006_/Q _4798_/Q _2779_/S vssd1 vssd1 vccd1 vccd1 _2777_/B sky130_fd_sc_hd__mux2_1
X_4446_ _4452_/A _4446_/B vssd1 vssd1 vccd1 vccd1 _4447_/A sky130_fd_sc_hd__and2_1
X_4377_ _4824_/Q _4812_/Q vssd1 vssd1 vccd1 vccd1 _4377_/Y sky130_fd_sc_hd__nand2_1
X_3328_ _3328_/A _3328_/B _3328_/C vssd1 vssd1 vccd1 vccd1 _3328_/X sky130_fd_sc_hd__and3_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _3241_/A _3245_/X _3248_/B _3256_/A _3246_/Y vssd1 vssd1 vccd1 vccd1 _3259_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_26_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5185__92 vssd1 vssd1 vccd1 vccd1 _5185__92/HI _5293_/A sky130_fd_sc_hd__conb_1
XFILLER_78_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2630_ _4964_/Q _4756_/Q _2639_/S vssd1 vssd1 vccd1 vccd1 _2631_/B sky130_fd_sc_hd__mux2_1
X_2561_ _4944_/Q _4736_/Q _2570_/S vssd1 vssd1 vccd1 vccd1 _2562_/B sky130_fd_sc_hd__mux2_1
X_2492_ _2516_/A vssd1 vssd1 vccd1 vccd1 _2497_/A sky130_fd_sc_hd__buf_6
X_5280_ _5280_/A _2475_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
X_4300_ _5013_/Q _4259_/X _4298_/Y _4299_/X _4281_/X vssd1 vssd1 vccd1 vccd1 _5013_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4231_ _4228_/X _4229_/Y _4230_/X vssd1 vssd1 vccd1 vccd1 _4231_/X sky130_fd_sc_hd__a21o_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4162_ _4996_/Q _4212_/B vssd1 vssd1 vccd1 vccd1 _4162_/X sky130_fd_sc_hd__or2_1
X_4093_ _4093_/A _4093_/B _4093_/C vssd1 vssd1 vccd1 vccd1 _4093_/X sky130_fd_sc_hd__and3_1
X_3113_ _4877_/Q _5045_/Q vssd1 vssd1 vccd1 vccd1 _3115_/A sky130_fd_sc_hd__or2_1
X_3044_ _4868_/Q _5036_/Q vssd1 vssd1 vccd1 vccd1 _3046_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4995_ _4995_/CLK _4995_/D vssd1 vssd1 vccd1 vccd1 _4995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3946_ _4969_/Q _3933_/X _3944_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _4969_/D sky130_fd_sc_hd__o211a_1
XFILLER_23_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3877_ _3842_/X _3874_/X _3875_/X _3876_/X vssd1 vssd1 vccd1 vccd1 _4960_/D sky130_fd_sc_hd__o211a_1
X_2828_ _2838_/A _2828_/B vssd1 vssd1 vccd1 vccd1 _2829_/A sky130_fd_sc_hd__and2_1
X_2759_ _5001_/Q _4793_/Q _2762_/S vssd1 vssd1 vccd1 vccd1 _2760_/B sky130_fd_sc_hd__mux2_1
X_4429_ _4435_/A _4429_/B vssd1 vssd1 vccd1 vccd1 _4430_/A sky130_fd_sc_hd__and2_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4780_ _4989_/CLK _4780_/D vssd1 vssd1 vccd1 vccd1 _4780_/Q sky130_fd_sc_hd__dfxtp_1
X_3800_ _4963_/Q _4743_/Q vssd1 vssd1 vccd1 vccd1 _3805_/C sky130_fd_sc_hd__or2_1
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3731_ _4941_/Q _3664_/A _3729_/Y _3730_/X _3646_/X vssd1 vssd1 vccd1 vccd1 _4941_/D
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_35_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5085_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3662_ _5113_/Q _4945_/Q vssd1 vssd1 vccd1 vccd1 _3663_/B sky130_fd_sc_hd__xnor2_1
X_2613_ _4959_/Q _4751_/Q _2622_/S vssd1 vssd1 vccd1 vccd1 _2614_/B sky130_fd_sc_hd__mux2_1
X_3593_ _3639_/B vssd1 vssd1 vccd1 vccd1 _3593_/X sky130_fd_sc_hd__clkbuf_2
X_2544_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2544_/Y sky130_fd_sc_hd__inv_2
X_2475_ _2478_/A vssd1 vssd1 vccd1 vccd1 _2475_/Y sky130_fd_sc_hd__inv_2
X_5263_ _5263_/A _2453_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
X_4214_ _4196_/A _4198_/Y _4203_/B _4211_/A _4201_/Y vssd1 vssd1 vccd1 vccd1 _4214_/Y
+ sky130_fd_sc_hd__a311oi_2
X_4145_ _4146_/A _4146_/B vssd1 vssd1 vccd1 vccd1 _4145_/X sky130_fd_sc_hd__or2_1
XFILLER_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4076_ _4076_/A vssd1 vssd1 vccd1 vccd1 _4076_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3027_ _4864_/Q _5032_/Q vssd1 vssd1 vccd1 vccd1 _3027_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4978_ _4978_/CLK _4978_/D vssd1 vssd1 vccd1 vccd1 _4978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3929_ _3921_/B _3926_/Y _3927_/Y _3878_/X vssd1 vssd1 vccd1 vccd1 _3929_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5155__62 vssd1 vssd1 vccd1 vccd1 _5155__62/HI _5250_/A sky130_fd_sc_hd__conb_1
XFILLER_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4901_ _5079_/CLK _4901_/D vssd1 vssd1 vccd1 vccd1 _4901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4832_ _4836_/CLK _4832_/D vssd1 vssd1 vccd1 vccd1 _5273_/A sky130_fd_sc_hd__dfxtp_1
X_4763_ _4981_/CLK _4763_/D vssd1 vssd1 vccd1 vccd1 _4763_/Q sky130_fd_sc_hd__dfxtp_1
X_4694_ _4694_/A vssd1 vssd1 vccd1 vccd1 _5110_/D sky130_fd_sc_hd__clkbuf_1
X_3714_ _3713_/Y _3695_/B _3693_/Y vssd1 vssd1 vccd1 vccd1 _3714_/Y sky130_fd_sc_hd__a21oi_1
X_3645_ _4022_/A vssd1 vssd1 vccd1 vccd1 _4076_/A sky130_fd_sc_hd__clkbuf_2
X_3576_ _3574_/X _3575_/Y _3558_/X vssd1 vssd1 vccd1 vccd1 _3576_/Y sky130_fd_sc_hd__a21oi_1
X_5315_ _5315_/A _2517_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2527_ _2527_/A vssd1 vssd1 vccd1 vccd1 _2527_/Y sky130_fd_sc_hd__inv_2
X_2458_ _2459_/A vssd1 vssd1 vccd1 vccd1 _2458_/Y sky130_fd_sc_hd__inv_2
X_5246_ _5246_/A _2545_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
X_4128_ _5004_/Q _4784_/Q vssd1 vssd1 vccd1 vccd1 _4135_/A sky130_fd_sc_hd__nand2_1
X_4059_ _4049_/A _4051_/Y _4057_/Y _4052_/X vssd1 vssd1 vccd1 vccd1 _4059_/X sky130_fd_sc_hd__a31o_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3430_ _3430_/A _3430_/B vssd1 vssd1 vccd1 vccd1 _3432_/B sky130_fd_sc_hd__and2_1
X_3361_ _3355_/Y _3272_/X _3358_/X _3359_/Y _3360_/X vssd1 vssd1 vccd1 vccd1 _4895_/D
+ sky130_fd_sc_hd__a221oi_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5103_/CLK _5100_/D vssd1 vssd1 vccd1 vccd1 _5100_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _4899_/Q _5067_/Q vssd1 vssd1 vccd1 vccd1 _3293_/B sky130_fd_sc_hd__and2_1
X_5031_ _5032_/CLK _5031_/D vssd1 vssd1 vccd1 vccd1 _5031_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5030_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4815_ _5027_/CLK _4815_/D vssd1 vssd1 vccd1 vccd1 _4815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4746_ _5122_/CLK _4746_/D vssd1 vssd1 vccd1 vccd1 _4746_/Q sky130_fd_sc_hd__dfxtp_1
X_4677_ _4677_/A vssd1 vssd1 vccd1 vccd1 _5105_/D sky130_fd_sc_hd__clkbuf_1
X_3628_ _4941_/Q _5109_/Q vssd1 vssd1 vccd1 vccd1 _3628_/Y sky130_fd_sc_hd__nor2_1
X_5125__32 vssd1 vssd1 vccd1 vccd1 _5125__32/HI _5220_/A sky130_fd_sc_hd__conb_1
X_3559_ _3555_/X _3563_/A _3558_/X vssd1 vssd1 vccd1 vccd1 _3559_/X sky130_fd_sc_hd__a21o_1
X_5229_ _5229_/A _2432_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2930_ _5277_/A _4852_/Q _2944_/S vssd1 vssd1 vccd1 vccd1 _2931_/B sky130_fd_sc_hd__mux2_1
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _4609_/A _4600_/B vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__and2_1
X_2861_ _2855_/X _4820_/Q _2557_/A _2860_/X vssd1 vssd1 vccd1 vccd1 _4820_/D sky130_fd_sc_hd__o211a_1
X_2792_ _5010_/Q _4802_/Q _2798_/S vssd1 vssd1 vccd1 vccd1 _2793_/B sky130_fd_sc_hd__mux2_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4531_ _4531_/A vssd1 vssd1 vccd1 vccd1 _5063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4462_ _4462_/A vssd1 vssd1 vccd1 vccd1 _5043_/D sky130_fd_sc_hd__clkbuf_1
X_3413_ _3411_/Y _3412_/X _3373_/X vssd1 vssd1 vccd1 vccd1 _3413_/X sky130_fd_sc_hd__a21o_1
X_4393_ _4384_/A _4386_/Y _4391_/X _4326_/X vssd1 vssd1 vccd1 vccd1 _4393_/X sky130_fd_sc_hd__a31o_1
X_3344_ _3336_/A _3338_/Y _3343_/X vssd1 vssd1 vccd1 vccd1 _3344_/Y sky130_fd_sc_hd__a21oi_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _4897_/Q _5065_/Q vssd1 vssd1 vccd1 vccd1 _3276_/B sky130_fd_sc_hd__xnor2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5015_/CLK _5014_/D vssd1 vssd1 vccd1 vccd1 _5014_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4729_ _4941_/Q _5121_/Q _4732_/S vssd1 vssd1 vccd1 vccd1 _4730_/B sky130_fd_sc_hd__mux2_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3060_ _3046_/A _3048_/Y _3053_/B _3051_/Y vssd1 vssd1 vccd1 vccd1 _3061_/B sky130_fd_sc_hd__a31o_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3962_ _4076_/A vssd1 vssd1 vccd1 vccd1 _3962_/X sky130_fd_sc_hd__buf_2
X_3893_ _3889_/X _3892_/X _3848_/X vssd1 vssd1 vccd1 vccd1 _3893_/X sky130_fd_sc_hd__a21o_1
X_2913_ _4030_/B _3168_/B _2965_/B vssd1 vssd1 vccd1 vccd1 _2967_/B sky130_fd_sc_hd__and3_1
X_2844_ _5025_/Q _4817_/Q _2850_/S vssd1 vssd1 vccd1 vccd1 _2845_/B sky130_fd_sc_hd__mux2_1
X_4514_ _4514_/A vssd1 vssd1 vccd1 vccd1 _5058_/D sky130_fd_sc_hd__clkbuf_1
X_2775_ _2775_/A vssd1 vssd1 vccd1 vccd1 _4797_/D sky130_fd_sc_hd__clkbuf_1
X_4445_ _4859_/Q _5039_/Q _4455_/S vssd1 vssd1 vccd1 vccd1 _4446_/B sky130_fd_sc_hd__mux2_1
X_4376_ _4376_/A _4376_/B _4376_/C vssd1 vssd1 vccd1 vccd1 _4376_/X sky130_fd_sc_hd__and3_1
X_3327_ _3327_/A _3327_/B _3331_/C vssd1 vssd1 vccd1 vccd1 _3328_/C sky130_fd_sc_hd__and3_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3258_ _3176_/X _3256_/X _3257_/X _3209_/X vssd1 vssd1 vccd1 vccd1 _4882_/D sky130_fd_sc_hd__o211a_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _3189_/A _3189_/B vssd1 vssd1 vccd1 vccd1 _3191_/B sky130_fd_sc_hd__and2_1
XFILLER_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2560_ _4281_/A vssd1 vssd1 vccd1 vccd1 _2575_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2491_ input1/X vssd1 vssd1 vccd1 vccd1 _2516_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _4230_/A vssd1 vssd1 vccd1 vccd1 _4230_/X sky130_fd_sc_hd__clkbuf_2
X_4161_ _4190_/A _4161_/B vssd1 vssd1 vccd1 vccd1 _4161_/X sky130_fd_sc_hd__xor2_1
XFILLER_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4092_ _4092_/A _4092_/B _4096_/C vssd1 vssd1 vccd1 vccd1 _4093_/C sky130_fd_sc_hd__and3_1
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3112_ _3138_/A _3109_/B _3105_/A vssd1 vssd1 vccd1 vccd1 _3116_/A sky130_fd_sc_hd__a21oi_1
X_3043_ _3013_/B _3040_/X _3042_/X vssd1 vssd1 vccd1 vccd1 _3048_/A sky130_fd_sc_hd__a21o_1
XFILLER_48_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _4995_/CLK _4994_/D vssd1 vssd1 vccd1 vccd1 _4994_/Q sky130_fd_sc_hd__dfxtp_1
X_3945_ _3945_/A vssd1 vssd1 vccd1 vccd1 _3945_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3876_ _3945_/A vssd1 vssd1 vccd1 vccd1 _3876_/X sky130_fd_sc_hd__clkbuf_2
X_2827_ _5020_/Q _4812_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _2828_/B sky130_fd_sc_hd__mux2_1
X_2758_ _2758_/A vssd1 vssd1 vccd1 vccd1 _4792_/D sky130_fd_sc_hd__clkbuf_1
X_2689_ _2696_/A _2689_/B vssd1 vssd1 vccd1 vccd1 _2690_/A sky130_fd_sc_hd__and2_1
X_4428_ _4854_/Q _5034_/Q _4438_/S vssd1 vssd1 vccd1 vccd1 _4429_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4359_ _5021_/Q _4400_/B vssd1 vssd1 vccd1 vccd1 _4359_/X sky130_fd_sc_hd__or2_1
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5027_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3730_ _3720_/A _3722_/Y _3728_/X _3680_/X vssd1 vssd1 vccd1 vccd1 _3730_/X sky130_fd_sc_hd__a31o_1
XFILLER_60_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3661_ _3737_/B vssd1 vssd1 vccd1 vccd1 _3664_/A sky130_fd_sc_hd__clkbuf_2
X_2612_ _2681_/A vssd1 vssd1 vccd1 vccd1 _2627_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3592_ _3558_/X _3590_/X _3591_/X _3566_/X vssd1 vssd1 vccd1 vccd1 _4924_/D sky130_fd_sc_hd__o211a_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2543_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2543_/Y sky130_fd_sc_hd__inv_2
X_5262_ _5262_/A _2452_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
X_2474_ _2478_/A vssd1 vssd1 vccd1 vccd1 _2474_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4213_ _4130_/X _4211_/X _4212_/X _4163_/X vssd1 vssd1 vccd1 vccd1 _5002_/D sky130_fd_sc_hd__o211a_1
X_4144_ _4144_/A _4144_/B vssd1 vssd1 vccd1 vccd1 _4146_/B sky130_fd_sc_hd__and2_1
XFILLER_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4075_ _4074_/A _4093_/B _4052_/X vssd1 vssd1 vccd1 vccd1 _4075_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3026_ _3020_/A _3019_/B _3024_/Y _3025_/Y vssd1 vssd1 vccd1 vccd1 _3026_/X sky130_fd_sc_hd__a211o_1
XFILLER_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4977_ _4978_/CLK _4977_/D vssd1 vssd1 vccd1 vccd1 _4977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3928_ _3921_/B _3926_/Y _3927_/Y vssd1 vssd1 vccd1 vccd1 _3928_/X sky130_fd_sc_hd__o21a_1
X_3859_ _3857_/X _3858_/Y _3842_/X vssd1 vssd1 vccd1 vccd1 _3859_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5170__77 vssd1 vssd1 vccd1 vccd1 _5170__77/HI _5265_/A sky130_fd_sc_hd__conb_1
XFILLER_59_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4900_ _5079_/CLK _4900_/D vssd1 vssd1 vccd1 vccd1 _4900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4831_ _5027_/CLK _4831_/D vssd1 vssd1 vccd1 vccd1 _4831_/Q sky130_fd_sc_hd__dfxtp_1
X_4762_ _4966_/CLK _4762_/D vssd1 vssd1 vccd1 vccd1 _4762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4693_ _4696_/A _4693_/B vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__and2_1
X_3713_ _5116_/Q _4948_/Q vssd1 vssd1 vccd1 vccd1 _3713_/Y sky130_fd_sc_hd__nand2_1
X_3644_ _3636_/B _3641_/Y _3642_/Y _3593_/X vssd1 vssd1 vccd1 vccd1 _3644_/Y sky130_fd_sc_hd__o31ai_1
X_3575_ _3575_/A _3575_/B vssd1 vssd1 vccd1 vccd1 _3575_/Y sky130_fd_sc_hd__nand2_1
X_5314_ _5314_/A _2515_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
X_2526_ _2527_/A vssd1 vssd1 vccd1 vccd1 _2526_/Y sky130_fd_sc_hd__inv_2
X_5245_ _5245_/A _2544_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_29_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2457_ _2459_/A vssd1 vssd1 vccd1 vccd1 _2457_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4127_ _5004_/Q _4784_/Q vssd1 vssd1 vccd1 vccd1 _4127_/X sky130_fd_sc_hd__or2_1
XFILLER_56_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4058_ _4049_/A _4051_/Y _4057_/Y vssd1 vssd1 vccd1 vccd1 _4058_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3009_ _3009_/A _3009_/B vssd1 vssd1 vccd1 vccd1 _3040_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3360_ _5285_/A vssd1 vssd1 vccd1 vccd1 _3360_/X sky130_fd_sc_hd__buf_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _4899_/Q _5067_/Q vssd1 vssd1 vccd1 vccd1 _3293_/A sky130_fd_sc_hd__nor2_1
X_5030_ _5030_/CLK _5030_/D vssd1 vssd1 vccd1 vccd1 _5030_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4814_ _5019_/CLK _4814_/D vssd1 vssd1 vccd1 vccd1 _4814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4745_ _4978_/CLK _4745_/D vssd1 vssd1 vccd1 vccd1 _4745_/Q sky130_fd_sc_hd__dfxtp_1
X_4676_ _4679_/A _4676_/B vssd1 vssd1 vccd1 vccd1 _4677_/A sky130_fd_sc_hd__and2_1
X_3627_ _4928_/Q _3554_/X _3626_/X _3566_/X vssd1 vssd1 vccd1 vccd1 _4928_/D sky130_fd_sc_hd__o211a_1
X_3558_ _3564_/A vssd1 vssd1 vccd1 vccd1 _3558_/X sky130_fd_sc_hd__clkbuf_2
X_2509_ _2509_/A vssd1 vssd1 vccd1 vccd1 _2509_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3489_ _3489_/A _3489_/B vssd1 vssd1 vccd1 vccd1 _3494_/A sky130_fd_sc_hd__nor2_1
X_5140__47 vssd1 vssd1 vccd1 vccd1 _5140__47/HI _5235_/A sky130_fd_sc_hd__conb_1
X_5228_ _5228_/A _2431_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2860_ _2858_/X _2859_/X _2855_/A vssd1 vssd1 vccd1 vccd1 _2860_/X sky130_fd_sc_hd__a21bo_1
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2791_ _2791_/A vssd1 vssd1 vccd1 vccd1 _4801_/D sky130_fd_sc_hd__clkbuf_1
X_4530_ _4539_/A _4530_/B vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__and2_1
X_4461_ _4470_/A _4461_/B vssd1 vssd1 vccd1 vccd1 _4462_/A sky130_fd_sc_hd__and2_1
X_3412_ _3421_/A _3412_/B vssd1 vssd1 vccd1 vccd1 _3412_/X sky130_fd_sc_hd__or2_1
X_4392_ _4384_/A _4386_/Y _4391_/X vssd1 vssd1 vccd1 vccd1 _4392_/Y sky130_fd_sc_hd__a21oi_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3341_/Y _3343_/B vssd1 vssd1 vccd1 vccd1 _3343_/X sky130_fd_sc_hd__and2b_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _4884_/Q _3268_/X _3273_/X _3209_/X vssd1 vssd1 vccd1 vccd1 _4884_/D sky130_fd_sc_hd__o211a_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5015_/CLK _5013_/D vssd1 vssd1 vccd1 vccd1 _5013_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2989_ _2986_/X _2987_/Y _2988_/X vssd1 vssd1 vccd1 vccd1 _2989_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4728_ _4728_/A vssd1 vssd1 vccd1 vccd1 _5120_/D sky130_fd_sc_hd__clkbuf_1
X_4659_ _4662_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4660_/A sky130_fd_sc_hd__and2_1
XFILLER_72_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5215__122 vssd1 vssd1 vccd1 vccd1 _5215__122/HI _5323_/A sky130_fd_sc_hd__conb_1
XFILLER_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5106_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ _3952_/A _3954_/Y _3959_/Y _3943_/X vssd1 vssd1 vccd1 vccd1 _3961_/X sky130_fd_sc_hd__a31o_1
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2912_ _3168_/A _4844_/Q vssd1 vssd1 vccd1 vccd1 _2965_/B sky130_fd_sc_hd__and2b_1
X_3892_ _3902_/A _3874_/B _3882_/A _3901_/A _3891_/Y vssd1 vssd1 vccd1 vccd1 _3892_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2843_ _2843_/A vssd1 vssd1 vccd1 vccd1 _4816_/D sky130_fd_sc_hd__clkbuf_1
X_2774_ _2784_/A _2774_/B vssd1 vssd1 vccd1 vccd1 _2775_/A sky130_fd_sc_hd__and2_1
X_4513_ _4522_/A _4513_/B vssd1 vssd1 vccd1 vccd1 _4514_/A sky130_fd_sc_hd__and2_1
X_4444_ _4444_/A vssd1 vssd1 vccd1 vccd1 _5038_/D sky130_fd_sc_hd__clkbuf_1
X_4375_ _4375_/A _4375_/B _4375_/C _4379_/C vssd1 vssd1 vccd1 vccd1 _4376_/C sky130_fd_sc_hd__and4_1
X_3326_ _4891_/Q _3277_/A _3323_/Y _3324_/X _3325_/X vssd1 vssd1 vccd1 vccd1 _4891_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _4882_/Q _3257_/B vssd1 vssd1 vccd1 vccd1 _3257_/X sky130_fd_sc_hd__or2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3188_ _4886_/Q _5054_/Q vssd1 vssd1 vccd1 vccd1 _3189_/B sky130_fd_sc_hd__or2_1
XFILLER_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5176__83 vssd1 vssd1 vccd1 vccd1 _5176__83/HI _5271_/A sky130_fd_sc_hd__conb_1
X_2490_ _2490_/A vssd1 vssd1 vccd1 vccd1 _2490_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ _4146_/A _4146_/B _4151_/Y _4159_/X vssd1 vssd1 vccd1 vccd1 _4161_/B sky130_fd_sc_hd__a31o_1
X_3111_ _3078_/X _3109_/X _3110_/X _3063_/X vssd1 vssd1 vccd1 vccd1 _4864_/D sky130_fd_sc_hd__o211a_1
X_4091_ _3992_/A _4043_/A _4089_/Y _4090_/X _4076_/X vssd1 vssd1 vccd1 vccd1 _4987_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3042_ _4867_/Q _5035_/Q _3028_/Y _3040_/C _3041_/X vssd1 vssd1 vccd1 vccd1 _3042_/X
+ sky130_fd_sc_hd__a221o_1
X_4993_ _4995_/CLK _4993_/D vssd1 vssd1 vccd1 vccd1 _4993_/Q sky130_fd_sc_hd__dfxtp_1
X_3944_ _3941_/X _3942_/Y _3943_/X vssd1 vssd1 vccd1 vccd1 _3944_/X sky130_fd_sc_hd__a21o_1
X_3875_ _4960_/Q _3924_/B vssd1 vssd1 vccd1 vccd1 _3875_/X sky130_fd_sc_hd__or2_1
X_2826_ _2826_/A vssd1 vssd1 vccd1 vccd1 _4811_/D sky130_fd_sc_hd__clkbuf_1
X_2757_ _2767_/A _2757_/B vssd1 vssd1 vccd1 vccd1 _2758_/A sky130_fd_sc_hd__and2_1
X_2688_ _4981_/Q _4773_/Q _2691_/S vssd1 vssd1 vccd1 vccd1 _2689_/B sky130_fd_sc_hd__mux2_1
X_4427_ _4427_/A vssd1 vssd1 vccd1 vccd1 _5033_/D sky130_fd_sc_hd__clkbuf_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _4358_/A _4376_/B vssd1 vssd1 vccd1 vccd1 _4358_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _3307_/Y _3309_/B vssd1 vssd1 vccd1 vccd1 _3328_/B sky130_fd_sc_hd__and2b_1
X_4289_ _5024_/Q _4804_/Q vssd1 vssd1 vccd1 vccd1 _4290_/B sky130_fd_sc_hd__or2_1
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ _4932_/Q _3652_/X _3657_/X _3659_/X vssd1 vssd1 vccd1 vccd1 _4932_/D sky130_fd_sc_hd__o211a_1
X_2611_ _2982_/A vssd1 vssd1 vccd1 vccd1 _2681_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3591_ _4924_/Q _3639_/B vssd1 vssd1 vccd1 vccd1 _3591_/X sky130_fd_sc_hd__or2_1
X_2542_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2542_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5261_ _5261_/A _2451_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
X_4212_ _5002_/Q _4212_/B vssd1 vssd1 vccd1 vccd1 _4212_/X sky130_fd_sc_hd__or2_1
X_2473_ _2485_/A vssd1 vssd1 vccd1 vccd1 _2478_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_44_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5058_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4143_ _5006_/Q _4786_/Q vssd1 vssd1 vccd1 vccd1 _4144_/B sky130_fd_sc_hd__or2_1
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4074_ _4074_/A _4093_/B vssd1 vssd1 vccd1 vccd1 _4074_/Y sky130_fd_sc_hd__nor2_1
X_3025_ _4865_/Q _5033_/Q vssd1 vssd1 vccd1 vccd1 _3025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4976_ _4978_/CLK _4976_/D vssd1 vssd1 vccd1 vccd1 _4976_/Q sky130_fd_sc_hd__dfxtp_1
X_3927_ _4979_/Q _4759_/Q vssd1 vssd1 vccd1 vccd1 _3927_/Y sky130_fd_sc_hd__xnor2_1
X_3858_ _3858_/A _3858_/B vssd1 vssd1 vccd1 vccd1 _3858_/Y sky130_fd_sc_hd__nand2_1
X_2809_ _5015_/Q _4807_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _2810_/B sky130_fd_sc_hd__mux2_1
X_3789_ _3789_/A _3806_/B vssd1 vssd1 vccd1 vccd1 _3789_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5146__53 vssd1 vssd1 vccd1 vccd1 _5146__53/HI _5241_/A sky130_fd_sc_hd__conb_1
XFILLER_41_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4830_ _4836_/CLK _4830_/D vssd1 vssd1 vccd1 vccd1 _4830_/Q sky130_fd_sc_hd__dfxtp_1
X_4761_ _4972_/CLK _4761_/D vssd1 vssd1 vccd1 vccd1 _4761_/Q sky130_fd_sc_hd__dfxtp_1
X_4692_ _4930_/Q _5110_/Q _4699_/S vssd1 vssd1 vccd1 vccd1 _4693_/B sky130_fd_sc_hd__mux2_1
X_3712_ _3712_/A _3712_/B _3712_/C vssd1 vssd1 vccd1 vccd1 _3712_/X sky130_fd_sc_hd__and3_1
X_3643_ _3636_/B _3641_/Y _3642_/Y vssd1 vssd1 vccd1 vccd1 _3643_/X sky130_fd_sc_hd__o21a_1
X_5313_ _5313_/A _2514_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
X_3574_ _3575_/A _3575_/B vssd1 vssd1 vccd1 vccd1 _3574_/X sky130_fd_sc_hd__or2_1
X_2525_ _2527_/A vssd1 vssd1 vccd1 vccd1 _2525_/Y sky130_fd_sc_hd__inv_2
X_2456_ _2459_/A vssd1 vssd1 vccd1 vccd1 _2456_/Y sky130_fd_sc_hd__inv_2
X_5244_ _5244_/A _2543_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
X_4126_ _4212_/B vssd1 vssd1 vccd1 vccd1 _4126_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4057_ _4057_/A _4057_/B vssd1 vssd1 vccd1 vccd1 _4057_/Y sky130_fd_sc_hd__nor2_1
X_3008_ _4864_/Q _5032_/Q vssd1 vssd1 vccd1 vccd1 _3009_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4959_ _4964_/CLK _4959_/D vssd1 vssd1 vccd1 vccd1 _4959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _4886_/Q _3268_/X _3289_/X _3279_/X vssd1 vssd1 vccd1 vccd1 _4886_/D sky130_fd_sc_hd__o211a_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4813_ _5050_/CLK _4813_/D vssd1 vssd1 vccd1 vccd1 _4813_/Q sky130_fd_sc_hd__dfxtp_1
X_4744_ _4978_/CLK _4744_/D vssd1 vssd1 vccd1 vccd1 _4744_/Q sky130_fd_sc_hd__dfxtp_1
X_4675_ _4925_/Q _5105_/Q _4682_/S vssd1 vssd1 vccd1 vccd1 _4676_/B sky130_fd_sc_hd__mux2_1
X_3626_ _3624_/X _3625_/Y _3564_/X vssd1 vssd1 vccd1 vccd1 _3626_/X sky130_fd_sc_hd__a21o_1
X_3557_ _3936_/A _3557_/B vssd1 vssd1 vccd1 vccd1 _3564_/A sky130_fd_sc_hd__or2_2
X_2508_ _2509_/A vssd1 vssd1 vccd1 vccd1 _2508_/Y sky130_fd_sc_hd__inv_2
X_5227_ _5227_/A _2428_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
X_3488_ _4924_/Q _5092_/Q vssd1 vssd1 vccd1 vccd1 _3489_/B sky130_fd_sc_hd__nor2_1
X_2439_ _2441_/A vssd1 vssd1 vccd1 vccd1 _2439_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4109_ _4101_/A _4103_/Y _4108_/X vssd1 vssd1 vccd1 vccd1 _4109_/Y sky130_fd_sc_hd__a21oi_1
X_5089_ _5091_/CLK _5089_/D vssd1 vssd1 vccd1 vccd1 _5089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2790_ _2803_/A _2790_/B vssd1 vssd1 vccd1 vccd1 _2791_/A sky130_fd_sc_hd__and2_1
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _4863_/Q _5043_/Q _4474_/S vssd1 vssd1 vccd1 vccd1 _4461_/B sky130_fd_sc_hd__mux2_1
X_3411_ _3421_/A _3412_/B vssd1 vssd1 vccd1 vccd1 _3411_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4391_ _4389_/Y _4391_/B vssd1 vssd1 vccd1 vccd1 _4391_/X sky130_fd_sc_hd__and2b_1
X_3342_ _4905_/Q _5073_/Q vssd1 vssd1 vccd1 vccd1 _3343_/B sky130_fd_sc_hd__nand2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3269_/X _3276_/A _3272_/X vssd1 vssd1 vccd1 vccd1 _3273_/X sky130_fd_sc_hd__a21o_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5015_/CLK _5012_/D vssd1 vssd1 vccd1 vccd1 _5012_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2988_ _2988_/A vssd1 vssd1 vccd1 vccd1 _2988_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4727_ _4730_/A _4727_/B vssd1 vssd1 vccd1 vccd1 _4728_/A sky130_fd_sc_hd__and2_1
X_4658_ _4920_/Q _5100_/Q _4665_/S vssd1 vssd1 vccd1 vccd1 _4659_/B sky130_fd_sc_hd__mux2_1
X_3609_ _4926_/Q _3554_/X _3608_/X _3566_/X vssd1 vssd1 vccd1 vccd1 _4926_/D sky130_fd_sc_hd__o211a_1
X_4589_ _4592_/A _4589_/B vssd1 vssd1 vccd1 vccd1 _4590_/A sky130_fd_sc_hd__and2_1
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3960_ _3952_/A _3954_/Y _3959_/Y vssd1 vssd1 vccd1 vccd1 _3960_/Y sky130_fd_sc_hd__a21oi_1
X_2911_ _4845_/Q vssd1 vssd1 vccd1 vccd1 _3168_/B sky130_fd_sc_hd__clkbuf_1
X_3891_ _3890_/Y _3882_/B _3888_/Y vssd1 vssd1 vccd1 vccd1 _3891_/Y sky130_fd_sc_hd__a21oi_1
X_2842_ _2917_/A _2842_/B vssd1 vssd1 vccd1 vccd1 _2843_/A sky130_fd_sc_hd__and2_1
X_2773_ _5005_/Q _4797_/Q _2779_/S vssd1 vssd1 vccd1 vccd1 _2774_/B sky130_fd_sc_hd__mux2_1
X_4512_ _4878_/Q _5058_/Q _4525_/S vssd1 vssd1 vccd1 vccd1 _4513_/B sky130_fd_sc_hd__mux2_1
X_4443_ _4452_/A _4443_/B vssd1 vssd1 vccd1 vccd1 _4444_/A sky130_fd_sc_hd__and2_1
X_4374_ _5023_/Q _4367_/A _4372_/Y _4373_/X _4281_/X vssd1 vssd1 vccd1 vccd1 _5023_/D
+ sky130_fd_sc_hd__o221a_1
X_3325_ _3551_/A vssd1 vssd1 vccd1 vccd1 _3325_/X sky130_fd_sc_hd__buf_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3256_/A _3256_/B vssd1 vssd1 vccd1 vccd1 _3256_/X sky130_fd_sc_hd__xor2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _4886_/Q _5054_/Q vssd1 vssd1 vccd1 vccd1 _3189_/A sky130_fd_sc_hd__nand2_1
X_5197__104 vssd1 vssd1 vccd1 vccd1 _5197__104/HI _5305_/A sky130_fd_sc_hd__conb_1
XFILLER_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5191__98 vssd1 vssd1 vccd1 vccd1 _5191__98/HI _5299_/A sky130_fd_sc_hd__conb_1
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3110_ _4864_/Q _3161_/B vssd1 vssd1 vccd1 vccd1 _3110_/X sky130_fd_sc_hd__or2_1
X_4090_ _4084_/Y _4086_/X _4092_/B _4096_/C _4052_/A vssd1 vssd1 vccd1 vccd1 _4090_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3041_ _4866_/Q _5034_/Q _3041_/C vssd1 vssd1 vccd1 vccd1 _3041_/X sky130_fd_sc_hd__and3_1
X_4992_ _4995_/CLK _4992_/D vssd1 vssd1 vccd1 vccd1 _4992_/Q sky130_fd_sc_hd__dfxtp_1
X_3943_ _3943_/A vssd1 vssd1 vccd1 vccd1 _3943_/X sky130_fd_sc_hd__clkbuf_2
X_3874_ _3902_/A _3874_/B vssd1 vssd1 vccd1 vccd1 _3874_/X sky130_fd_sc_hd__xor2_1
XFILLER_31_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2825_ _2838_/A _2825_/B vssd1 vssd1 vccd1 vccd1 _2826_/A sky130_fd_sc_hd__and2_1
X_2756_ _5000_/Q _4792_/Q _2762_/S vssd1 vssd1 vccd1 vccd1 _2757_/B sky130_fd_sc_hd__mux2_1
X_2687_ _2687_/A vssd1 vssd1 vccd1 vccd1 _4772_/D sky130_fd_sc_hd__clkbuf_1
X_4426_ _4435_/A _4426_/B vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__and2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _4355_/Y _4357_/B vssd1 vssd1 vccd1 vccd1 _4376_/B sky130_fd_sc_hd__and2b_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _4901_/Q _5069_/Q vssd1 vssd1 vccd1 vccd1 _3309_/B sky130_fd_sc_hd__nand2_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _5024_/Q _4804_/Q vssd1 vssd1 vccd1 vccd1 _4290_/A sky130_fd_sc_hd__nand2_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _4892_/Q _5060_/Q vssd1 vssd1 vccd1 vccd1 _3241_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2610_ _2610_/A vssd1 vssd1 vccd1 vccd1 _4750_/D sky130_fd_sc_hd__clkbuf_1
X_3590_ _3617_/A _3590_/B vssd1 vssd1 vccd1 vccd1 _3590_/X sky130_fd_sc_hd__xor2_1
X_2541_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2541_/Y sky130_fd_sc_hd__inv_2
X_2472_ _2472_/A vssd1 vssd1 vccd1 vccd1 _2472_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5260_ _5260_/A _2450_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4211_ _4211_/A _4211_/B vssd1 vssd1 vccd1 vccd1 _4211_/X sky130_fd_sc_hd__xor2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4142_ _5006_/Q _4786_/Q vssd1 vssd1 vccd1 vccd1 _4144_/A sky130_fd_sc_hd__nand2_1
X_4073_ _4071_/Y _4073_/B vssd1 vssd1 vccd1 vccd1 _4093_/B sky130_fd_sc_hd__and2b_1
X_3024_ _3039_/A vssd1 vssd1 vccd1 vccd1 _3024_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5004_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4975_ _4975_/CLK _4975_/D vssd1 vssd1 vccd1 vccd1 _4975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3926_ _3908_/A _3910_/Y _3915_/B _3923_/A _3913_/Y vssd1 vssd1 vccd1 vccd1 _3926_/Y
+ sky130_fd_sc_hd__a311oi_2
X_3857_ _3858_/A _3858_/B vssd1 vssd1 vccd1 vccd1 _3857_/X sky130_fd_sc_hd__or2_1
X_2808_ _2808_/A vssd1 vssd1 vccd1 vccd1 _4806_/D sky130_fd_sc_hd__clkbuf_1
X_3788_ _3786_/Y _3788_/B vssd1 vssd1 vccd1 vccd1 _3806_/B sky130_fd_sc_hd__and2b_1
X_2739_ _4995_/Q _4787_/Q _2745_/S vssd1 vssd1 vccd1 vccd1 _2740_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4409_ _4418_/A _4409_/B vssd1 vssd1 vccd1 vccd1 _4410_/A sky130_fd_sc_hd__and2_1
XFILLER_74_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5161__68 vssd1 vssd1 vccd1 vccd1 _5161__68/HI _5256_/A sky130_fd_sc_hd__conb_1
XFILLER_73_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4760_ _4978_/CLK _4760_/D vssd1 vssd1 vccd1 vccd1 _4760_/Q sky130_fd_sc_hd__dfxtp_1
X_4691_ _4691_/A vssd1 vssd1 vccd1 vccd1 _5109_/D sky130_fd_sc_hd__clkbuf_1
X_3711_ _3711_/A _3711_/B _3711_/C vssd1 vssd1 vccd1 vccd1 _3712_/C sky130_fd_sc_hd__and3_1
X_3642_ _5111_/Q _4943_/Q vssd1 vssd1 vccd1 vccd1 _3642_/Y sky130_fd_sc_hd__xnor2_1
X_5312_ _5312_/A _2513_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
X_3573_ _3573_/A _3573_/B vssd1 vssd1 vccd1 vccd1 _3575_/B sky130_fd_sc_hd__and2_1
X_2524_ _2527_/A vssd1 vssd1 vccd1 vccd1 _2524_/Y sky130_fd_sc_hd__inv_2
X_2455_ _2459_/A vssd1 vssd1 vccd1 vccd1 _2455_/Y sky130_fd_sc_hd__inv_2
X_5243_ _5243_/A _2542_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_68_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4125_ _4125_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _4212_/B sky130_fd_sc_hd__nor2_2
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4056_ _4995_/Q _4775_/Q vssd1 vssd1 vccd1 vccd1 _4057_/B sky130_fd_sc_hd__and2_1
X_3007_ _4864_/Q _5032_/Q vssd1 vssd1 vccd1 vccd1 _3009_/A sky130_fd_sc_hd__and2_1
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _4964_/CLK _4958_/D vssd1 vssd1 vccd1 vccd1 _4958_/Q sky130_fd_sc_hd__dfxtp_1
X_3909_ _3910_/A _3910_/B vssd1 vssd1 vccd1 vccd1 _3909_/X sky130_fd_sc_hd__or2_1
X_4889_ _5070_/CLK _4889_/D vssd1 vssd1 vccd1 vccd1 _4889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4812_ _5019_/CLK _4812_/D vssd1 vssd1 vccd1 vccd1 _4812_/Q sky130_fd_sc_hd__dfxtp_1
X_4743_ _4954_/CLK _4743_/D vssd1 vssd1 vccd1 vccd1 _4743_/Q sky130_fd_sc_hd__dfxtp_1
X_4674_ _4674_/A vssd1 vssd1 vccd1 vccd1 _5104_/D sky130_fd_sc_hd__clkbuf_1
X_3625_ _3625_/A _3625_/B vssd1 vssd1 vccd1 vccd1 _3625_/Y sky130_fd_sc_hd__nand2_2
X_3556_ _4932_/Q _5100_/Q vssd1 vssd1 vccd1 vccd1 _3563_/A sky130_fd_sc_hd__nand2_1
X_2507_ _2509_/A vssd1 vssd1 vccd1 vccd1 _2507_/Y sky130_fd_sc_hd__inv_2
X_5226_ _5226_/A _2427_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
X_3487_ _4924_/Q _5092_/Q vssd1 vssd1 vccd1 vccd1 _3489_/A sky130_fd_sc_hd__and2_1
X_2438_ _2441_/A vssd1 vssd1 vccd1 vccd1 _2438_/Y sky130_fd_sc_hd__inv_2
X_4108_ _4106_/Y _4108_/B vssd1 vssd1 vccd1 vccd1 _4108_/X sky130_fd_sc_hd__and2b_1
X_5088_ _5091_/CLK _5088_/D vssd1 vssd1 vccd1 vccd1 _5088_/Q sky130_fd_sc_hd__dfxtp_1
X_4039_ _4035_/X _4042_/A _4038_/X vssd1 vssd1 vccd1 vccd1 _4039_/X sky130_fd_sc_hd__a21o_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5131__38 vssd1 vssd1 vccd1 vccd1 _5131__38/HI _5226_/A sky130_fd_sc_hd__conb_1
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3410_ _3406_/A _3405_/B _3403_/Y vssd1 vssd1 vccd1 vccd1 _3412_/B sky130_fd_sc_hd__a21oi_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4390_ _4829_/Q _4817_/Q vssd1 vssd1 vccd1 vccd1 _4391_/B sky130_fd_sc_hd__nand2_1
X_3341_ _4905_/Q _5073_/Q vssd1 vssd1 vccd1 vccd1 _3341_/Y sky130_fd_sc_hd__nor2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _3288_/A vssd1 vssd1 vccd1 vccd1 _3272_/X sky130_fd_sc_hd__clkbuf_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5011_ _5026_/CLK _5011_/D vssd1 vssd1 vccd1 vccd1 _5011_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2987_ _2987_/A _2987_/B vssd1 vssd1 vccd1 vccd1 _2987_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4726_ _4940_/Q _5120_/Q _4732_/S vssd1 vssd1 vccd1 vccd1 _4727_/B sky130_fd_sc_hd__mux2_1
X_4657_ _4657_/A vssd1 vssd1 vccd1 vccd1 _5099_/D sky130_fd_sc_hd__clkbuf_1
X_3608_ _3604_/X _3607_/X _3564_/X vssd1 vssd1 vccd1 vccd1 _3608_/X sky130_fd_sc_hd__a21o_1
X_4588_ _4900_/Q _5080_/Q _4595_/S vssd1 vssd1 vccd1 vccd1 _4589_/B sky130_fd_sc_hd__mux2_1
X_3539_ _4930_/Q _5098_/Q vssd1 vssd1 vccd1 vccd1 _3541_/A sky130_fd_sc_hd__or2_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2910_ _4846_/Q vssd1 vssd1 vccd1 vccd1 _4030_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3890_ _4972_/Q _4752_/Q vssd1 vssd1 vccd1 vccd1 _3890_/Y sky130_fd_sc_hd__nand2_1
X_2841_ _5024_/Q _4816_/Q _2850_/S vssd1 vssd1 vccd1 vccd1 _2842_/B sky130_fd_sc_hd__mux2_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2772_ _2772_/A vssd1 vssd1 vccd1 vccd1 _4796_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5087_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4511_ _4528_/A vssd1 vssd1 vccd1 vccd1 _4525_/S sky130_fd_sc_hd__buf_2
XFILLER_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4442_ _4858_/Q _5038_/Q _4455_/S vssd1 vssd1 vccd1 vccd1 _4443_/B sky130_fd_sc_hd__mux2_1
X_4373_ _4375_/B _4369_/X _4375_/C _4379_/C _4326_/X vssd1 vssd1 vccd1 vccd1 _4373_/X
+ sky130_fd_sc_hd__a41o_1
X_3324_ _3318_/Y _3320_/X _3327_/B _3331_/C _3288_/A vssd1 vssd1 vccd1 vccd1 _3324_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3241_/A _3245_/X _3248_/B _3246_/Y vssd1 vssd1 vccd1 vccd1 _3256_/B sky130_fd_sc_hd__a31o_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3181_/A _3181_/B _3185_/Y vssd1 vssd1 vccd1 vccd1 _3191_/A sky130_fd_sc_hd__o21ai_1
XFILLER_26_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_4709_ _4935_/Q _5115_/Q _4716_/S vssd1 vssd1 vccd1 vccd1 _4710_/B sky130_fd_sc_hd__mux2_1
XFILLER_1_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3040_ _3040_/A _3040_/B _3040_/C vssd1 vssd1 vccd1 vccd1 _3040_/X sky130_fd_sc_hd__and3_1
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _5018_/CLK _4991_/D vssd1 vssd1 vccd1 vccd1 _4991_/Q sky130_fd_sc_hd__dfxtp_1
X_3942_ _3942_/A _3942_/B vssd1 vssd1 vccd1 vccd1 _3942_/Y sky130_fd_sc_hd__nand2_1
X_3873_ _3858_/A _3858_/B _3863_/Y _3872_/X vssd1 vssd1 vccd1 vccd1 _3874_/B sky130_fd_sc_hd__a31o_1
X_2824_ _5019_/Q _4811_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _2825_/B sky130_fd_sc_hd__mux2_1
X_2755_ _2755_/A vssd1 vssd1 vccd1 vccd1 _4791_/D sky130_fd_sc_hd__clkbuf_1
X_5167__74 vssd1 vssd1 vccd1 vccd1 _5167__74/HI _5262_/A sky130_fd_sc_hd__conb_1
XFILLER_8_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2686_ _2696_/A _2686_/B vssd1 vssd1 vccd1 vccd1 _2687_/A sky130_fd_sc_hd__and2_1
X_4425_ _4853_/Q _5033_/Q _4438_/S vssd1 vssd1 vccd1 vccd1 _4426_/B sky130_fd_sc_hd__mux2_1
X_4356_ _4825_/Q _4813_/Q vssd1 vssd1 vccd1 vccd1 _4357_/B sky130_fd_sc_hd__nand2_1
X_3307_ _4901_/Q _5069_/Q vssd1 vssd1 vccd1 vccd1 _3307_/Y sky130_fd_sc_hd__nor2_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5205__112 vssd1 vssd1 vccd1 vccd1 _5205__112/HI _5313_/A sky130_fd_sc_hd__conb_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _4256_/B _4284_/X _4286_/X vssd1 vssd1 vccd1 vccd1 _4292_/A sky130_fd_sc_hd__a21o_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _3207_/B _3233_/X _3237_/X vssd1 vssd1 vccd1 vccd1 _3242_/A sky130_fd_sc_hd__a21o_1
X_3169_ _3936_/A vssd1 vssd1 vccd1 vccd1 _4318_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2540_ _2540_/A vssd1 vssd1 vccd1 vccd1 _2545_/A sky130_fd_sc_hd__buf_8
X_2471_ _2472_/A vssd1 vssd1 vccd1 vccd1 _2471_/Y sky130_fd_sc_hd__inv_2
X_4210_ _4196_/A _4198_/Y _4203_/B _4201_/Y vssd1 vssd1 vccd1 vccd1 _4211_/B sky130_fd_sc_hd__a31o_1
X_4141_ _4135_/A _4135_/B _4140_/Y vssd1 vssd1 vccd1 vccd1 _4146_/A sky130_fd_sc_hd__o21ai_1
X_4072_ _4997_/Q _4777_/Q vssd1 vssd1 vccd1 vccd1 _4073_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3023_ _4866_/Q _5034_/Q vssd1 vssd1 vccd1 vccd1 _3039_/A sky130_fd_sc_hd__xor2_1
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4974_ _4981_/CLK _4974_/D vssd1 vssd1 vccd1 vccd1 _4974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3925_ _3842_/X _3923_/X _3924_/X _3876_/X vssd1 vssd1 vccd1 vccd1 _4966_/D sky130_fd_sc_hd__o211a_1
X_3856_ _3856_/A _3856_/B vssd1 vssd1 vccd1 vccd1 _3858_/B sky130_fd_sc_hd__and2_1
X_3787_ _4961_/Q _4741_/Q vssd1 vssd1 vccd1 vccd1 _3788_/B sky130_fd_sc_hd__nand2_1
X_2807_ _2821_/A _2807_/B vssd1 vssd1 vccd1 vccd1 _2808_/A sky130_fd_sc_hd__and2_1
X_2738_ _2738_/A vssd1 vssd1 vccd1 vccd1 _4786_/D sky130_fd_sc_hd__clkbuf_1
X_2669_ _2679_/A _2669_/B vssd1 vssd1 vccd1 vccd1 _2670_/A sky130_fd_sc_hd__and2_1
X_4408_ _4848_/Q _5028_/Q _4421_/S vssd1 vssd1 vccd1 vccd1 _4409_/B sky130_fd_sc_hd__mux2_1
X_4339_ _4823_/Q _4811_/Q vssd1 vssd1 vccd1 vccd1 _4341_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3710_ _4939_/Q _3664_/A _3708_/Y _3709_/X _3646_/X vssd1 vssd1 vccd1 vccd1 _4939_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4690_ _4696_/A _4690_/B vssd1 vssd1 vccd1 vccd1 _4691_/A sky130_fd_sc_hd__and2_1
X_3641_ _3623_/A _3625_/Y _3630_/B _3638_/A _3628_/Y vssd1 vssd1 vccd1 vccd1 _3641_/Y
+ sky130_fd_sc_hd__a311oi_2
X_3572_ _4934_/Q _5102_/Q vssd1 vssd1 vccd1 vccd1 _3573_/B sky130_fd_sc_hd__or2_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5137__44 vssd1 vssd1 vccd1 vccd1 _5137__44/HI _5232_/A sky130_fd_sc_hd__conb_1
X_5311_ _5311_/A _2512_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
X_2523_ _2527_/A vssd1 vssd1 vccd1 vccd1 _2523_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5242_ _5242_/A _2541_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
X_2454_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2459_/A sky130_fd_sc_hd__buf_8
XFILLER_68_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4124_ _4119_/Y _4038_/X _4122_/X _4123_/Y _3360_/X vssd1 vssd1 vccd1 vccd1 _4991_/D
+ sky130_fd_sc_hd__a221oi_1
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4055_ _4995_/Q _4775_/Q vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3006_ _4851_/Q _2976_/X _3004_/Y _3005_/X _2897_/X vssd1 vssd1 vccd1 vccd1 _4851_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4957_ _4964_/CLK _4957_/D vssd1 vssd1 vccd1 vccd1 _4957_/Q sky130_fd_sc_hd__dfxtp_1
X_3908_ _3908_/A _3908_/B vssd1 vssd1 vccd1 vccd1 _3910_/B sky130_fd_sc_hd__and2_1
X_4888_ _5070_/CLK _4888_/D vssd1 vssd1 vccd1 vccd1 _4888_/Q sky130_fd_sc_hd__dfxtp_1
X_3839_ _4968_/Q _4748_/Q vssd1 vssd1 vccd1 vccd1 _3839_/X sky130_fd_sc_hd__or2_1
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4811_ _5019_/CLK _4811_/D vssd1 vssd1 vccd1 vccd1 _4811_/Q sky130_fd_sc_hd__dfxtp_1
X_4742_ _4954_/CLK _4742_/D vssd1 vssd1 vccd1 vccd1 _4742_/Q sky130_fd_sc_hd__dfxtp_1
X_4673_ _4679_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4674_/A sky130_fd_sc_hd__and2_1
X_3624_ _3625_/A _3625_/B vssd1 vssd1 vccd1 vccd1 _3624_/X sky130_fd_sc_hd__or2_1
X_3555_ _4932_/Q _5100_/Q vssd1 vssd1 vccd1 vccd1 _3555_/X sky130_fd_sc_hd__or2_1
X_2506_ _2509_/A vssd1 vssd1 vccd1 vccd1 _2506_/Y sky130_fd_sc_hd__inv_2
X_3486_ _4911_/Q _3457_/A _3484_/Y _3485_/X _3441_/X vssd1 vssd1 vccd1 vccd1 _4911_/D
+ sky130_fd_sc_hd__o221a_1
X_2437_ _2441_/A vssd1 vssd1 vccd1 vccd1 _2437_/Y sky130_fd_sc_hd__inv_2
X_5225_ _5225_/A _2426_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4107_ _5001_/Q _4781_/Q vssd1 vssd1 vccd1 vccd1 _4108_/B sky130_fd_sc_hd__nand2_1
X_5087_ _5087_/CLK _5087_/D vssd1 vssd1 vccd1 vccd1 _5087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4038_ _4052_/A vssd1 vssd1 vccd1 vccd1 _4038_/X sky130_fd_sc_hd__clkbuf_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3340_ _4892_/Q _3268_/X _3339_/X _3279_/X vssd1 vssd1 vccd1 vccd1 _4892_/D sky130_fd_sc_hd__o211a_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _4037_/A _3553_/B vssd1 vssd1 vccd1 vccd1 _3288_/A sky130_fd_sc_hd__or2_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5010_/CLK _5010_/D vssd1 vssd1 vccd1 vccd1 _5010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2986_ _2987_/A _2987_/B vssd1 vssd1 vccd1 vccd1 _2986_/X sky130_fd_sc_hd__or2_1
X_4725_ _4725_/A vssd1 vssd1 vccd1 vccd1 _5119_/D sky130_fd_sc_hd__clkbuf_1
X_4656_ _4662_/A _4656_/B vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__and2_1
X_4587_ _4587_/A vssd1 vssd1 vccd1 vccd1 _5079_/D sky130_fd_sc_hd__clkbuf_1
X_3607_ _3617_/A _3590_/B _3597_/A _3616_/A _3606_/Y vssd1 vssd1 vccd1 vccd1 _3607_/X
+ sky130_fd_sc_hd__a311o_1
X_3538_ _4917_/Q _3457_/A _3536_/Y _3537_/X _3441_/X vssd1 vssd1 vccd1 vccd1 _4917_/D
+ sky130_fd_sc_hd__o221a_1
X_3469_ _4909_/Q _3457_/X _3468_/X _3434_/X vssd1 vssd1 vccd1 vccd1 _4909_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_8_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4999_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2840_ _2919_/A vssd1 vssd1 vccd1 vccd1 _2917_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2771_ _2784_/A _2771_/B vssd1 vssd1 vccd1 vccd1 _2772_/A sky130_fd_sc_hd__and2_1
X_4510_ _4510_/A vssd1 vssd1 vccd1 vccd1 _5057_/D sky130_fd_sc_hd__clkbuf_1
X_4441_ _4441_/A vssd1 vssd1 vccd1 vccd1 _4455_/S sky130_fd_sc_hd__buf_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ _4375_/B _4369_/X _4375_/C _4379_/C vssd1 vssd1 vccd1 vccd1 _4372_/Y sky130_fd_sc_hd__a22oi_1
X_3323_ _3318_/Y _3320_/X _3327_/B _3331_/C vssd1 vssd1 vccd1 vccd1 _3323_/Y sky130_fd_sc_hd__a22oi_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _3254_/A _3254_/B vssd1 vssd1 vccd1 vccd1 _3256_/A sky130_fd_sc_hd__nand2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _4885_/Q _5053_/Q vssd1 vssd1 vccd1 vccd1 _3185_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2969_ _3648_/A _2967_/B _2968_/Y vssd1 vssd1 vccd1 vccd1 _4847_/D sky130_fd_sc_hd__o21a_1
X_4708_ _4708_/A vssd1 vssd1 vccd1 vccd1 _5114_/D sky130_fd_sc_hd__clkbuf_1
X_4639_ _4639_/A vssd1 vssd1 vccd1 vccd1 _5094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _5018_/CLK _4990_/D vssd1 vssd1 vccd1 vccd1 _4990_/Q sky130_fd_sc_hd__dfxtp_1
X_3941_ _3942_/A _3942_/B vssd1 vssd1 vccd1 vccd1 _3941_/X sky130_fd_sc_hd__or2_1
X_3872_ _4970_/Q _4750_/Q _3871_/X _3863_/B vssd1 vssd1 vccd1 vccd1 _3872_/X sky130_fd_sc_hd__a31o_1
XFILLER_31_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2823_ _2919_/A vssd1 vssd1 vccd1 vccd1 _2838_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2754_ _2767_/A _2754_/B vssd1 vssd1 vccd1 vccd1 _2755_/A sky130_fd_sc_hd__and2_1
X_2685_ _4980_/Q _4772_/Q _2691_/S vssd1 vssd1 vccd1 vccd1 _2686_/B sky130_fd_sc_hd__mux2_1
X_4424_ _4441_/A vssd1 vssd1 vccd1 vccd1 _4438_/S sky130_fd_sc_hd__buf_2
X_5182__89 vssd1 vssd1 vccd1 vccd1 _5182__89/HI _5290_/A sky130_fd_sc_hd__conb_1
X_4355_ _4825_/Q _4813_/Q vssd1 vssd1 vccd1 vccd1 _4355_/Y sky130_fd_sc_hd__nor2_1
X_3306_ _3328_/A _3303_/B _3299_/A vssd1 vssd1 vccd1 vccd1 _3310_/A sky130_fd_sc_hd__a21oi_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _5023_/Q _4803_/Q _4272_/Y _4284_/C _4285_/X vssd1 vssd1 vccd1 vccd1 _4286_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _4891_/Q _5059_/Q _3235_/Y _3233_/C _3236_/X vssd1 vssd1 vccd1 vccd1 _3237_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3168_ _3168_/A _3168_/B _4844_/Q vssd1 vssd1 vccd1 vccd1 _3936_/A sky130_fd_sc_hd__or3_2
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3099_ _3099_/A _3099_/B vssd1 vssd1 vccd1 vccd1 _3099_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2470_ _2472_/A vssd1 vssd1 vccd1 vccd1 _2470_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4140_ _5005_/Q _4785_/Q vssd1 vssd1 vccd1 vccd1 _4140_/Y sky130_fd_sc_hd__nand2_1
X_4071_ _4997_/Q _4777_/Q vssd1 vssd1 vccd1 vccd1 _4071_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3022_ _4853_/Q _2976_/A _3020_/Y _3021_/X _2897_/X vssd1 vssd1 vccd1 vccd1 _4853_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _4981_/CLK _4973_/D vssd1 vssd1 vccd1 vccd1 _4973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3924_ _4966_/Q _3924_/B vssd1 vssd1 vccd1 vccd1 _3924_/X sky130_fd_sc_hd__or2_1
X_3855_ _4970_/Q _4750_/Q vssd1 vssd1 vccd1 vccd1 _3856_/B sky130_fd_sc_hd__or2_1
X_3786_ _4961_/Q _4741_/Q vssd1 vssd1 vccd1 vccd1 _3786_/Y sky130_fd_sc_hd__nor2_1
X_2806_ _5014_/Q _4806_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _2807_/B sky130_fd_sc_hd__mux2_1
X_2737_ _2750_/A _2737_/B vssd1 vssd1 vccd1 vccd1 _2738_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4964_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2668_ _4975_/Q _4767_/Q _2674_/S vssd1 vssd1 vccd1 vccd1 _2669_/B sky130_fd_sc_hd__mux2_1
X_4407_ _4441_/A vssd1 vssd1 vccd1 vccd1 _4421_/S sky130_fd_sc_hd__buf_2
X_2599_ _2609_/A _2599_/B vssd1 vssd1 vccd1 vccd1 _2600_/A sky130_fd_sc_hd__and2_1
X_4338_ _4319_/X _4336_/X _4337_/X _4321_/X vssd1 vssd1 vccd1 vccd1 _5018_/D sky130_fd_sc_hd__o211a_1
XFILLER_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4269_ _5021_/Q _4801_/Q vssd1 vssd1 vccd1 vccd1 _4269_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3640_ _3558_/X _3638_/X _3639_/X _3566_/X vssd1 vssd1 vccd1 vccd1 _4930_/D sky130_fd_sc_hd__o211a_1
X_3571_ _4934_/Q _5102_/Q vssd1 vssd1 vccd1 vccd1 _3573_/A sky130_fd_sc_hd__nand2_1
X_2522_ _2540_/A vssd1 vssd1 vccd1 vccd1 _2527_/A sky130_fd_sc_hd__buf_8
X_5310_ _5310_/A _2511_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5241_ _5241_/A _2539_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
X_2453_ _2453_/A vssd1 vssd1 vccd1 vccd1 _2453_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5152__59 vssd1 vssd1 vccd1 vccd1 _5152__59/HI _5247_/A sky130_fd_sc_hd__conb_1
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4123_ _4114_/B _4120_/X _4121_/X _4052_/X vssd1 vssd1 vccd1 vccd1 _4123_/Y sky130_fd_sc_hd__a31oi_1
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
X_4054_ _4982_/Q _4034_/X _4053_/X _4023_/X vssd1 vssd1 vccd1 vccd1 _4982_/D sky130_fd_sc_hd__o211a_1
X_3005_ _2996_/A _2998_/Y _3003_/Y _2988_/X vssd1 vssd1 vccd1 vccd1 _3005_/X sky130_fd_sc_hd__a31o_1
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ _4964_/CLK _4956_/D vssd1 vssd1 vccd1 vccd1 _4956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3907_ _4976_/Q _4756_/Q vssd1 vssd1 vccd1 vccd1 _3908_/B sky130_fd_sc_hd__or2_1
X_4887_ _5070_/CLK _4887_/D vssd1 vssd1 vccd1 vccd1 _4887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3838_ _3924_/B vssd1 vssd1 vccd1 vccd1 _3838_/X sky130_fd_sc_hd__clkbuf_2
X_3769_ _4959_/Q _4739_/Q vssd1 vssd1 vccd1 vccd1 _3770_/B sky130_fd_sc_hd__and2_1
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _5018_/CLK _4810_/D vssd1 vssd1 vccd1 vccd1 _4810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4741_ _4948_/CLK _4741_/D vssd1 vssd1 vccd1 vccd1 _4741_/Q sky130_fd_sc_hd__dfxtp_1
X_4672_ _4924_/Q _5104_/Q _4682_/S vssd1 vssd1 vccd1 vccd1 _4673_/B sky130_fd_sc_hd__mux2_1
X_3623_ _3623_/A _3623_/B vssd1 vssd1 vccd1 vccd1 _3625_/B sky130_fd_sc_hd__and2_1
X_3554_ _3639_/B vssd1 vssd1 vccd1 vccd1 _3554_/X sky130_fd_sc_hd__clkbuf_2
X_2505_ _2509_/A vssd1 vssd1 vccd1 vccd1 _2505_/Y sky130_fd_sc_hd__inv_2
X_3485_ _3475_/A _3477_/Y _3483_/Y _3467_/X vssd1 vssd1 vccd1 vccd1 _3485_/X sky130_fd_sc_hd__a31o_1
X_5224_ _5224_/A _2425_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
X_2436_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2441_/A sky130_fd_sc_hd__buf_12
X_4106_ _5001_/Q _4781_/Q vssd1 vssd1 vccd1 vccd1 _4106_/Y sky130_fd_sc_hd__nor2_1
X_5086_ _5087_/CLK _5086_/D vssd1 vssd1 vccd1 vccd1 _5086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4037_ _4037_/A _4223_/B vssd1 vssd1 vccd1 vccd1 _4052_/A sky130_fd_sc_hd__or2_2
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4939_ _4954_/CLK _4939_/D vssd1 vssd1 vccd1 vccd1 _4939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3270_ _4896_/Q _5064_/Q vssd1 vssd1 vccd1 vccd1 _3276_/A sky130_fd_sc_hd__nand2_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2985_ _4861_/Q _5029_/Q vssd1 vssd1 vccd1 vccd1 _2987_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4724_ _4730_/A _4724_/B vssd1 vssd1 vccd1 vccd1 _4725_/A sky130_fd_sc_hd__and2_1
X_4655_ _4919_/Q _5099_/Q _4665_/S vssd1 vssd1 vccd1 vccd1 _4656_/B sky130_fd_sc_hd__mux2_1
X_4586_ _4592_/A _4586_/B vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__and2_1
X_3606_ _3605_/Y _3597_/B _3603_/Y vssd1 vssd1 vccd1 vccd1 _3606_/Y sky130_fd_sc_hd__a21oi_1
X_3537_ _3528_/A _3530_/X _3535_/X _3467_/A vssd1 vssd1 vccd1 vccd1 _3537_/X sky130_fd_sc_hd__a31o_1
X_3468_ _3465_/X _3466_/Y _3467_/X vssd1 vssd1 vccd1 vccd1 _3468_/X sky130_fd_sc_hd__a21o_1
X_2419_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2419_/Y sky130_fd_sc_hd__inv_2
X_3399_ _4900_/Q _3448_/B vssd1 vssd1 vccd1 vccd1 _3399_/X sky130_fd_sc_hd__or2_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5069_ _5077_/CLK _5069_/D vssd1 vssd1 vccd1 vccd1 _5069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5188__95 vssd1 vssd1 vccd1 vccd1 _5188__95/HI _5296_/A sky130_fd_sc_hd__conb_1
XFILLER_4_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2770_ _5004_/Q _4796_/Q _2779_/S vssd1 vssd1 vccd1 vccd1 _2771_/B sky130_fd_sc_hd__mux2_1
X_4440_ _4440_/A vssd1 vssd1 vccd1 vccd1 _5037_/D sky130_fd_sc_hd__clkbuf_1
X_4371_ _4827_/Q _4815_/Q vssd1 vssd1 vccd1 vccd1 _4379_/C sky130_fd_sc_hd__or2_1
X_3322_ _4903_/Q _5071_/Q vssd1 vssd1 vccd1 vccd1 _3331_/C sky130_fd_sc_hd__or2_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _4894_/Q _5062_/Q vssd1 vssd1 vccd1 vccd1 _3254_/B sky130_fd_sc_hd__nand2_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5033_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3184_ _4873_/Q _3172_/X _3183_/X _3148_/X vssd1 vssd1 vccd1 vccd1 _4873_/D sky130_fd_sc_hd__o211a_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2968_ _5285_/A _2968_/B vssd1 vssd1 vccd1 vccd1 _2968_/Y sky130_fd_sc_hd__nor2_1
X_4707_ _4713_/A _4707_/B vssd1 vssd1 vccd1 vccd1 _4708_/A sky130_fd_sc_hd__and2_1
X_4638_ _4644_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _4639_/A sky130_fd_sc_hd__and2_1
X_2899_ _2886_/X input12/X _2887_/X vssd1 vssd1 vccd1 vccd1 _2899_/X sky130_fd_sc_hd__o21a_1
X_4569_ _4575_/A _4569_/B vssd1 vssd1 vccd1 vccd1 _4570_/A sky130_fd_sc_hd__and2_1
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _4981_/Q _4761_/Q vssd1 vssd1 vccd1 vccd1 _3942_/B sky130_fd_sc_hd__xnor2_1
XFILLER_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3871_ _4971_/Q _4751_/Q vssd1 vssd1 vccd1 vccd1 _3871_/X sky130_fd_sc_hd__or2_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2822_ _2822_/A vssd1 vssd1 vccd1 vccd1 _4810_/D sky130_fd_sc_hd__clkbuf_1
X_2753_ _4999_/Q _4791_/Q _2762_/S vssd1 vssd1 vccd1 vccd1 _2754_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2684_ _2684_/A vssd1 vssd1 vccd1 vccd1 _4771_/D sky130_fd_sc_hd__clkbuf_1
X_4423_ _4423_/A vssd1 vssd1 vccd1 vccd1 _5032_/D sky130_fd_sc_hd__clkbuf_1
X_4354_ _4376_/A _4351_/B _4347_/A vssd1 vssd1 vccd1 vccd1 _4358_/A sky130_fd_sc_hd__a21oi_1
X_3305_ _3272_/X _3303_/X _3304_/X _3279_/X vssd1 vssd1 vccd1 vccd1 _4888_/D sky130_fd_sc_hd__o211a_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _5022_/Q _4802_/Q _4285_/C vssd1 vssd1 vccd1 vccd1 _4285_/X sky130_fd_sc_hd__and3_1
XFILLER_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3236_ _4890_/Q _5058_/Q _3236_/C vssd1 vssd1 vccd1 vccd1 _3236_/X sky130_fd_sc_hd__and3_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3167_ _4871_/Q _3074_/A _3165_/Y _3166_/X _3135_/X vssd1 vssd1 vccd1 vccd1 _4871_/D
+ sky130_fd_sc_hd__o221a_1
X_3098_ _4875_/Q _5043_/Q vssd1 vssd1 vccd1 vccd1 _3099_/B sky130_fd_sc_hd__and2_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5158__65 vssd1 vssd1 vccd1 vccd1 _5158__65/HI _5253_/A sky130_fd_sc_hd__conb_1
XFILLER_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _4093_/A _4067_/B _4063_/A vssd1 vssd1 vccd1 vccd1 _4074_/A sky130_fd_sc_hd__a21oi_1
X_3021_ _3020_/A _3040_/B _2988_/X vssd1 vssd1 vccd1 vccd1 _3021_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4972_ _4972_/CLK _4972_/D vssd1 vssd1 vccd1 vccd1 _4972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3923_ _3923_/A _3923_/B vssd1 vssd1 vccd1 vccd1 _3923_/X sky130_fd_sc_hd__xor2_1
X_3854_ _4970_/Q _4750_/Q vssd1 vssd1 vccd1 vccd1 _3856_/A sky130_fd_sc_hd__nand2_1
X_2805_ _2919_/A vssd1 vssd1 vccd1 vccd1 _2821_/A sky130_fd_sc_hd__clkbuf_2
X_3785_ _3806_/A _3781_/B _3777_/A vssd1 vssd1 vccd1 vccd1 _3789_/A sky130_fd_sc_hd__a21oi_1
X_2736_ _4994_/Q _4786_/Q _2745_/S vssd1 vssd1 vccd1 vccd1 _2737_/B sky130_fd_sc_hd__mux2_1
X_2667_ _2667_/A vssd1 vssd1 vccd1 vccd1 _4766_/D sky130_fd_sc_hd__clkbuf_1
X_4406_ _5027_/Q _4367_/A _4404_/X _4405_/Y _2557_/A vssd1 vssd1 vccd1 vccd1 _5027_/D
+ sky130_fd_sc_hd__o221a_1
X_2598_ _4955_/Q _4747_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _2599_/B sky130_fd_sc_hd__mux2_1
X_4337_ _5018_/Q _4400_/B vssd1 vssd1 vccd1 vccd1 _4337_/X sky130_fd_sc_hd__or2_1
X_4268_ _4283_/A vssd1 vssd1 vccd1 vccd1 _4268_/Y sky130_fd_sc_hd__inv_2
X_3219_ _4890_/Q _5058_/Q vssd1 vssd1 vccd1 vccd1 _3232_/B sky130_fd_sc_hd__nand2_1
X_4199_ _4197_/X _4198_/Y _4136_/X vssd1 vssd1 vccd1 vccd1 _4199_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3570_ _3563_/A _3563_/B _3569_/Y vssd1 vssd1 vccd1 vccd1 _3575_/A sky130_fd_sc_hd__o21ai_1
X_2521_ _2521_/A vssd1 vssd1 vccd1 vccd1 _2521_/Y sky130_fd_sc_hd__inv_2
X_5240_ _5240_/A _2538_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2452_ _2453_/A vssd1 vssd1 vccd1 vccd1 _2452_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4114_/B _4120_/X _4121_/X vssd1 vssd1 vccd1 vccd1 _4122_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4053_ _4050_/X _4051_/Y _4052_/X vssd1 vssd1 vccd1 vccd1 _4053_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
X_3004_ _2996_/A _2998_/Y _3003_/Y vssd1 vssd1 vccd1 vccd1 _3004_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4955_ _5122_/CLK _4955_/D vssd1 vssd1 vccd1 vccd1 _4955_/Q sky130_fd_sc_hd__dfxtp_1
X_3906_ _4976_/Q _4756_/Q vssd1 vssd1 vccd1 vccd1 _3908_/A sky130_fd_sc_hd__nand2_1
X_4886_ _5070_/CLK _4886_/D vssd1 vssd1 vccd1 vccd1 _4886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3837_ _4219_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _3924_/B sky130_fd_sc_hd__nor2_2
X_3768_ _4959_/Q _4739_/Q vssd1 vssd1 vccd1 vccd1 _3770_/A sky130_fd_sc_hd__nor2_1
X_2719_ _2733_/A _2719_/B vssd1 vssd1 vccd1 vccd1 _2720_/A sky130_fd_sc_hd__and2_1
X_5128__35 vssd1 vssd1 vccd1 vccd1 _5128__35/HI _5223_/A sky130_fd_sc_hd__conb_1
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3699_ _5118_/Q _4950_/Q vssd1 vssd1 vccd1 vccd1 _3711_/A sky130_fd_sc_hd__xor2_1
XFILLER_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4740_ _4964_/CLK _4740_/D vssd1 vssd1 vccd1 vccd1 _4740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4671_ _4671_/A vssd1 vssd1 vccd1 vccd1 _5103_/D sky130_fd_sc_hd__clkbuf_1
X_3622_ _4940_/Q _5108_/Q vssd1 vssd1 vccd1 vccd1 _3623_/B sky130_fd_sc_hd__or2_1
X_3553_ _4318_/A _3553_/B vssd1 vssd1 vccd1 vccd1 _3639_/B sky130_fd_sc_hd__nor2_2
X_2504_ _2516_/A vssd1 vssd1 vccd1 vccd1 _2509_/A sky130_fd_sc_hd__buf_8
X_3484_ _3475_/A _3477_/Y _3483_/Y vssd1 vssd1 vccd1 vccd1 _3484_/Y sky130_fd_sc_hd__a21oi_1
X_2435_ _2435_/A vssd1 vssd1 vccd1 vccd1 _2435_/Y sky130_fd_sc_hd__inv_2
X_5223_ _5223_/A _2424_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
X_4105_ _4988_/Q _4034_/X _4104_/X _4082_/X vssd1 vssd1 vccd1 vccd1 _4988_/D sky130_fd_sc_hd__o211a_1
X_5085_ _5085_/CLK _5085_/D vssd1 vssd1 vccd1 vccd1 _5085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4036_ _4992_/Q _4772_/Q vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__nand2_1
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4938_ _4954_/CLK _4938_/D vssd1 vssd1 vccd1 vccd1 _4938_/Q sky130_fd_sc_hd__dfxtp_1
X_4869_ _5062_/CLK _4869_/D vssd1 vssd1 vccd1 vccd1 _4869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2984_ _4848_/Q _2976_/X _2981_/X _2983_/X vssd1 vssd1 vccd1 vccd1 _4848_/D sky130_fd_sc_hd__o211a_1
XFILLER_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4723_ _4939_/Q _5119_/Q _4732_/S vssd1 vssd1 vccd1 vccd1 _4724_/B sky130_fd_sc_hd__mux2_1
X_4654_ _4654_/A vssd1 vssd1 vccd1 vccd1 _5098_/D sky130_fd_sc_hd__clkbuf_1
X_4585_ _4899_/Q _5079_/Q _4595_/S vssd1 vssd1 vccd1 vccd1 _4586_/B sky130_fd_sc_hd__mux2_1
X_3605_ _4936_/Q _5104_/Q vssd1 vssd1 vccd1 vccd1 _3605_/Y sky130_fd_sc_hd__nand2_1
X_3536_ _3528_/A _3530_/X _3535_/X vssd1 vssd1 vccd1 vccd1 _3536_/Y sky130_fd_sc_hd__a21oi_1
X_3467_ _3467_/A vssd1 vssd1 vccd1 vccd1 _3467_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3398_ _3422_/A _3398_/B vssd1 vssd1 vccd1 vccd1 _3398_/X sky130_fd_sc_hd__xor2_1
X_2418_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2418_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5068_ _5077_/CLK _5068_/D vssd1 vssd1 vccd1 vccd1 _5068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4019_ _4005_/X _4018_/Y _4010_/A vssd1 vssd1 vccd1 vccd1 _4020_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4370_ _4827_/Q _4815_/Q vssd1 vssd1 vccd1 vccd1 _4375_/C sky130_fd_sc_hd__nand2_1
X_3321_ _4903_/Q _5071_/Q vssd1 vssd1 vccd1 vccd1 _3327_/B sky130_fd_sc_hd__nand2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3252_ _4894_/Q _5062_/Q vssd1 vssd1 vccd1 vccd1 _3254_/A sky130_fd_sc_hd__or2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _3180_/X _3181_/Y _3182_/X vssd1 vssd1 vccd1 vccd1 _3183_/X sky130_fd_sc_hd__a21o_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4978_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2967_ _2967_/A _2967_/B _2967_/C vssd1 vssd1 vccd1 vccd1 _4846_/D sky130_fd_sc_hd__nor3_1
X_2898_ _2878_/X _4828_/Q _2895_/X _2896_/X _2897_/X vssd1 vssd1 vccd1 vccd1 _4828_/D
+ sky130_fd_sc_hd__o221a_1
X_4706_ _4934_/Q _5114_/Q _4716_/S vssd1 vssd1 vccd1 vccd1 _4707_/B sky130_fd_sc_hd__mux2_1
X_4637_ _4914_/Q _5094_/Q _4648_/S vssd1 vssd1 vccd1 vccd1 _4638_/B sky130_fd_sc_hd__mux2_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4568_ _4894_/Q _5074_/Q _4578_/S vssd1 vssd1 vccd1 vccd1 _4569_/B sky130_fd_sc_hd__mux2_1
X_4499_ _4505_/A _4499_/B vssd1 vssd1 vccd1 vccd1 _4500_/A sky130_fd_sc_hd__and2_1
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3519_ _4915_/Q _3457_/A _3515_/X _3518_/X _3441_/X vssd1 vssd1 vccd1 vccd1 _4915_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ _3870_/A _3870_/B vssd1 vssd1 vccd1 vccd1 _3902_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2821_ _2821_/A _2821_/B vssd1 vssd1 vccd1 vccd1 _2822_/A sky130_fd_sc_hd__and2_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2752_ _2769_/A vssd1 vssd1 vccd1 vccd1 _2767_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4422_ _4435_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _4423_/A sky130_fd_sc_hd__and2_1
X_2683_ _2696_/A _2683_/B vssd1 vssd1 vccd1 vccd1 _2684_/A sky130_fd_sc_hd__and2_1
X_4353_ _4319_/X _4351_/X _4352_/X _4321_/X vssd1 vssd1 vccd1 vccd1 _5020_/D sky130_fd_sc_hd__o211a_1
X_3304_ _4888_/Q _3352_/B vssd1 vssd1 vccd1 vccd1 _3304_/X sky130_fd_sc_hd__or2_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4284_ _4284_/A _4284_/B _4284_/C vssd1 vssd1 vccd1 vccd1 _4284_/X sky130_fd_sc_hd__and3_1
X_3235_ _3234_/Y _3214_/B _3212_/Y vssd1 vssd1 vccd1 vccd1 _3235_/Y sky130_fd_sc_hd__a21oi_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3166_ _3158_/B _3163_/X _3164_/X _3084_/A vssd1 vssd1 vccd1 vccd1 _3166_/X sky130_fd_sc_hd__a31o_1
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3097_ _4875_/Q _5043_/Q vssd1 vssd1 vccd1 vccd1 _3099_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3999_ _3998_/Y _3976_/Y _3997_/B _3977_/A vssd1 vssd1 vccd1 vccd1 _3999_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5212__119 vssd1 vssd1 vccd1 vccd1 _5212__119/HI _5320_/A sky130_fd_sc_hd__conb_1
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3020_ _3020_/A _3040_/B vssd1 vssd1 vccd1 vccd1 _3020_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4971_ _4981_/CLK _4971_/D vssd1 vssd1 vccd1 vccd1 _4971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3922_ _3908_/A _3910_/Y _3915_/B _3913_/Y vssd1 vssd1 vccd1 vccd1 _3923_/B sky130_fd_sc_hd__a31o_1
X_3853_ _3847_/A _3847_/B _3852_/Y vssd1 vssd1 vccd1 vccd1 _3858_/A sky130_fd_sc_hd__o21ai_1
X_2804_ _2804_/A vssd1 vssd1 vccd1 vccd1 _4805_/D sky130_fd_sc_hd__clkbuf_1
X_3784_ _3830_/B vssd1 vssd1 vccd1 vccd1 _3784_/X sky130_fd_sc_hd__clkbuf_2
X_2735_ _2769_/A vssd1 vssd1 vccd1 vccd1 _2750_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2666_ _2679_/A _2666_/B vssd1 vssd1 vccd1 vccd1 _2667_/A sky130_fd_sc_hd__and2_1
X_4405_ _4397_/B _4402_/Y _4403_/Y _4367_/A vssd1 vssd1 vccd1 vccd1 _4405_/Y sky130_fd_sc_hd__o31ai_1
X_4336_ _4336_/A _4336_/B vssd1 vssd1 vccd1 vccd1 _4336_/X sky130_fd_sc_hd__and2_1
X_2597_ _2597_/A vssd1 vssd1 vccd1 vccd1 _4746_/D sky130_fd_sc_hd__clkbuf_1
X_4267_ _5022_/Q _4802_/Q vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__xor2_2
X_4198_ _4198_/A _4198_/B vssd1 vssd1 vccd1 vccd1 _4198_/Y sky130_fd_sc_hd__nand2_2
X_3218_ _4890_/Q _5058_/Q vssd1 vssd1 vccd1 vccd1 _3232_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5101_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3149_ _4868_/Q _3074_/X _3147_/X _3148_/X vssd1 vssd1 vccd1 vccd1 _4868_/D sky130_fd_sc_hd__o211a_1
XFILLER_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5193__100 vssd1 vssd1 vccd1 vccd1 _5193__100/HI _5301_/A sky130_fd_sc_hd__conb_1
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2520_ _2521_/A vssd1 vssd1 vccd1 vccd1 _2520_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2451_ _2453_/A vssd1 vssd1 vccd1 vccd1 _2451_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4121_ _5003_/Q _4783_/Q vssd1 vssd1 vccd1 vccd1 _4121_/X sky130_fd_sc_hd__xor2_1
X_4052_ _4052_/A vssd1 vssd1 vccd1 vccd1 _4052_/X sky130_fd_sc_hd__clkbuf_2
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
X_3003_ _3003_/A _3003_/B vssd1 vssd1 vccd1 vccd1 _3003_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4954_ _4954_/CLK _4954_/D vssd1 vssd1 vccd1 vccd1 _4954_/Q sky130_fd_sc_hd__dfxtp_1
X_3905_ _3874_/B _3902_/X _3904_/X vssd1 vssd1 vccd1 vccd1 _3910_/A sky130_fd_sc_hd__a21o_1
XFILLER_20_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4885_ _5070_/CLK _4885_/D vssd1 vssd1 vccd1 vccd1 _4885_/Q sky130_fd_sc_hd__dfxtp_1
X_3836_ _4955_/Q _3784_/X _3834_/X _3835_/Y _3773_/X vssd1 vssd1 vccd1 vccd1 _4955_/D
+ sky130_fd_sc_hd__o221a_1
X_3767_ _3758_/Y _3749_/X _3766_/Y _3479_/X vssd1 vssd1 vccd1 vccd1 _4946_/D sky130_fd_sc_hd__a211oi_1
X_2718_ _4989_/Q _4781_/Q _2727_/S vssd1 vssd1 vccd1 vccd1 _2719_/B sky130_fd_sc_hd__mux2_1
X_3698_ _4937_/Q _3652_/X _3697_/X _3659_/X vssd1 vssd1 vccd1 vccd1 _4937_/D sky130_fd_sc_hd__o211a_1
X_2649_ _2662_/A _2649_/B vssd1 vssd1 vccd1 vccd1 _2650_/A sky130_fd_sc_hd__and2_1
X_5299_ _5299_/A _2497_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
X_4319_ _4326_/A vssd1 vssd1 vccd1 vccd1 _4319_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _4679_/A _4670_/B vssd1 vssd1 vccd1 vccd1 _4671_/A sky130_fd_sc_hd__and2_1
X_3621_ _4940_/Q _5108_/Q vssd1 vssd1 vccd1 vccd1 _3623_/A sky130_fd_sc_hd__nand2_2
X_3552_ _4919_/Q _3457_/A _3549_/Y _3550_/X _3551_/X vssd1 vssd1 vccd1 vccd1 _4919_/D
+ sky130_fd_sc_hd__o221a_1
X_2503_ _2503_/A vssd1 vssd1 vccd1 vccd1 _2503_/Y sky130_fd_sc_hd__inv_2
X_3483_ _3483_/A _3483_/B vssd1 vssd1 vccd1 vccd1 _3483_/Y sky130_fd_sc_hd__nor2_1
X_2434_ _2435_/A vssd1 vssd1 vccd1 vccd1 _2434_/Y sky130_fd_sc_hd__inv_2
X_5222_ _5222_/A _2422_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
X_4104_ _4102_/X _4103_/Y _4052_/X vssd1 vssd1 vccd1 vccd1 _4104_/X sky130_fd_sc_hd__a21o_1
X_5084_ _5085_/CLK _5084_/D vssd1 vssd1 vccd1 vccd1 _5084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4035_ _4992_/Q _4772_/Q vssd1 vssd1 vccd1 vccd1 _4035_/X sky130_fd_sc_hd__or2_1
XFILLER_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4937_ _5117_/CLK _4937_/D vssd1 vssd1 vccd1 vccd1 _4937_/Q sky130_fd_sc_hd__dfxtp_1
X_4868_ _5048_/CLK _4868_/D vssd1 vssd1 vccd1 vccd1 _4868_/Q sky130_fd_sc_hd__dfxtp_1
X_3819_ _4965_/Q _4745_/Q vssd1 vssd1 vccd1 vccd1 _3819_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4799_ _5004_/CLK _4799_/D vssd1 vssd1 vccd1 vccd1 _4799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2983_ _4733_/A vssd1 vssd1 vccd1 vccd1 _2983_/X sky130_fd_sc_hd__clkbuf_2
X_4722_ _4722_/A vssd1 vssd1 vccd1 vccd1 _5118_/D sky130_fd_sc_hd__clkbuf_1
X_4653_ _4662_/A _4653_/B vssd1 vssd1 vccd1 vccd1 _4654_/A sky130_fd_sc_hd__and2_1
X_4584_ _4584_/A vssd1 vssd1 vccd1 vccd1 _5078_/D sky130_fd_sc_hd__clkbuf_1
X_3604_ _3598_/A _3597_/B _3602_/Y _3603_/Y vssd1 vssd1 vccd1 vccd1 _3604_/X sky130_fd_sc_hd__a211o_1
X_3535_ _3533_/Y _3535_/B vssd1 vssd1 vccd1 vccd1 _3535_/X sky130_fd_sc_hd__and2b_1
X_3466_ _3466_/A _3466_/B vssd1 vssd1 vccd1 vccd1 _3466_/Y sky130_fd_sc_hd__nand2_1
X_2417_ _2548_/A vssd1 vssd1 vccd1 vccd1 _2422_/A sky130_fd_sc_hd__buf_12
X_3397_ _3383_/A _3383_/B _3388_/Y _3396_/X vssd1 vssd1 vccd1 vccd1 _3398_/B sky130_fd_sc_hd__a31o_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5067_ _5077_/CLK _5067_/D vssd1 vssd1 vccd1 vccd1 _5067_/Q sky130_fd_sc_hd__dfxtp_1
X_4018_ _4988_/Q _4768_/Q _4010_/B vssd1 vssd1 vccd1 vccd1 _4018_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5179__86 vssd1 vssd1 vccd1 vccd1 _5179__86/HI _5287_/A sky130_fd_sc_hd__conb_1
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3320_ _3320_/A _3320_/B vssd1 vssd1 vccd1 vccd1 _3320_/X sky130_fd_sc_hd__or2_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _4881_/Q _3223_/A _3249_/Y _3250_/X _3230_/X vssd1 vssd1 vccd1 vccd1 _4881_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _3182_/A vssd1 vssd1 vccd1 vccd1 _3182_/X sky130_fd_sc_hd__buf_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2966_ _4030_/B _2966_/B vssd1 vssd1 vccd1 vccd1 _2967_/C sky130_fd_sc_hd__nor2_1
X_2897_ _3037_/A vssd1 vssd1 vccd1 vccd1 _2897_/X sky130_fd_sc_hd__buf_2
X_4705_ _4705_/A vssd1 vssd1 vccd1 vccd1 _5113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4636_ _4636_/A vssd1 vssd1 vccd1 vccd1 _5093_/D sky130_fd_sc_hd__clkbuf_1
X_4567_ _4567_/A vssd1 vssd1 vccd1 vccd1 _5073_/D sky130_fd_sc_hd__clkbuf_1
X_4498_ _4874_/Q _5054_/Q _4508_/S vssd1 vssd1 vccd1 vccd1 _4499_/B sky130_fd_sc_hd__mux2_1
X_3518_ _3520_/A _3507_/X _3516_/Y _3517_/X _3467_/A vssd1 vssd1 vccd1 vccd1 _3518_/X
+ sky130_fd_sc_hd__a41o_1
X_3449_ _3367_/X _3447_/X _3448_/X _3434_/X vssd1 vssd1 vccd1 vccd1 _4906_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5119_ _5121_/CLK _5119_/D vssd1 vssd1 vccd1 vccd1 _5119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2820_ _5018_/Q _4810_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _2821_/B sky130_fd_sc_hd__mux2_1
X_2751_ _2751_/A vssd1 vssd1 vccd1 vccd1 _4790_/D sky130_fd_sc_hd__clkbuf_1
X_2682_ _4979_/Q _4771_/Q _2691_/S vssd1 vssd1 vccd1 vccd1 _2683_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4421_ _4852_/Q _5032_/Q _4421_/S vssd1 vssd1 vccd1 vccd1 _4422_/B sky130_fd_sc_hd__mux2_1
X_4352_ _5020_/Q _4400_/B vssd1 vssd1 vccd1 vccd1 _4352_/X sky130_fd_sc_hd__or2_1
X_3303_ _3328_/A _3303_/B vssd1 vssd1 vccd1 vccd1 _3303_/X sky130_fd_sc_hd__xor2_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4283_ _4283_/A _4283_/B _4285_/C vssd1 vssd1 vccd1 vccd1 _4284_/C sky130_fd_sc_hd__and3_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _4888_/Q _5056_/Q vssd1 vssd1 vccd1 vccd1 _3234_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3165_ _3158_/B _3163_/X _3164_/X vssd1 vssd1 vccd1 vccd1 _3165_/Y sky130_fd_sc_hd__a21oi_1
X_3096_ _3087_/Y _3078_/X _3095_/Y _2967_/A vssd1 vssd1 vccd1 vccd1 _4862_/D sky130_fd_sc_hd__a211oi_1
XFILLER_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3998_ _4984_/Q _4764_/Q vssd1 vssd1 vccd1 vccd1 _3998_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2949_ _2949_/A vssd1 vssd1 vccd1 vccd1 _4841_/D sky130_fd_sc_hd__clkbuf_1
X_4619_ _4909_/Q _5089_/Q _4629_/S vssd1 vssd1 vccd1 vccd1 _4620_/B sky130_fd_sc_hd__mux2_1
XFILLER_77_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5149__56 vssd1 vssd1 vccd1 vccd1 _5149__56/HI _5244_/A sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_1_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5040_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _4972_/CLK _4970_/D vssd1 vssd1 vccd1 vccd1 _4970_/Q sky130_fd_sc_hd__dfxtp_1
X_3921_ _3921_/A _3921_/B vssd1 vssd1 vccd1 vccd1 _3923_/A sky130_fd_sc_hd__or2_1
X_3852_ _4969_/Q _4749_/Q vssd1 vssd1 vccd1 vccd1 _3852_/Y sky130_fd_sc_hd__nand2_1
X_2803_ _2803_/A _2803_/B vssd1 vssd1 vccd1 vccd1 _2804_/A sky130_fd_sc_hd__and2_1
X_3783_ _3749_/X _3781_/X _3782_/X _3724_/X vssd1 vssd1 vccd1 vccd1 _4948_/D sky130_fd_sc_hd__o211a_1
X_2734_ _2734_/A vssd1 vssd1 vccd1 vccd1 _4785_/D sky130_fd_sc_hd__clkbuf_1
X_2665_ _4974_/Q _4766_/Q _2674_/S vssd1 vssd1 vccd1 vccd1 _2666_/B sky130_fd_sc_hd__mux2_1
X_4404_ _4397_/B _4402_/Y _4403_/Y vssd1 vssd1 vccd1 vccd1 _4404_/X sky130_fd_sc_hd__o21a_1
X_2596_ _2609_/A _2596_/B vssd1 vssd1 vccd1 vccd1 _2597_/A sky130_fd_sc_hd__and2_1
X_5163__70 vssd1 vssd1 vccd1 vccd1 _5163__70/HI _5258_/A sky130_fd_sc_hd__conb_1
X_4335_ _4335_/A _4335_/B vssd1 vssd1 vccd1 vccd1 _4336_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4266_ _5009_/Q _4259_/X _4264_/Y _4265_/X _4187_/X vssd1 vssd1 vccd1 vccd1 _5009_/D
+ sky130_fd_sc_hd__o221a_1
X_4197_ _4198_/A _4198_/B vssd1 vssd1 vccd1 vccd1 _4197_/X sky130_fd_sc_hd__or2_1
X_3217_ _4877_/Q _3172_/X _3215_/Y _3216_/X _3135_/X vssd1 vssd1 vccd1 vccd1 _4877_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3148_ _4733_/A vssd1 vssd1 vccd1 vccd1 _3148_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3079_ _3075_/X _3083_/A _3078_/X vssd1 vssd1 vccd1 vccd1 _3079_/X sky130_fd_sc_hd__a21o_1
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2450_ _2453_/A vssd1 vssd1 vccd1 vccd1 _2450_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4120_ _4101_/A _4103_/Y _4108_/B _4116_/A _4106_/Y vssd1 vssd1 vccd1 vccd1 _4120_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_83_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ _4051_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _4051_/Y sky130_fd_sc_hd__nand2_1
X_3002_ _4863_/Q _5031_/Q vssd1 vssd1 vccd1 vccd1 _3003_/B sky130_fd_sc_hd__and2_1
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4953_ _4978_/CLK _4953_/D vssd1 vssd1 vccd1 vccd1 _4953_/Q sky130_fd_sc_hd__dfxtp_1
X_3904_ _4975_/Q _4755_/Q _3891_/Y _3902_/C _3903_/X vssd1 vssd1 vccd1 vccd1 _3904_/X
+ sky130_fd_sc_hd__a221o_1
X_4884_ _5070_/CLK _4884_/D vssd1 vssd1 vccd1 vccd1 _4884_/Q sky130_fd_sc_hd__dfxtp_1
X_3835_ _3827_/B _3832_/Y _3833_/Y _3784_/X vssd1 vssd1 vccd1 vccd1 _3835_/Y sky130_fd_sc_hd__o31ai_1
X_3766_ _3764_/X _3765_/Y _3749_/X vssd1 vssd1 vccd1 vccd1 _3766_/Y sky130_fd_sc_hd__a21oi_1
X_2717_ _2769_/A vssd1 vssd1 vccd1 vccd1 _2733_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3697_ _3692_/Y _3712_/B _3696_/Y vssd1 vssd1 vccd1 vccd1 _3697_/X sky130_fd_sc_hd__a21o_1
X_2648_ _4969_/Q _4761_/Q _2657_/S vssd1 vssd1 vccd1 vccd1 _2649_/B sky130_fd_sc_hd__mux2_1
X_2579_ _2592_/A _2579_/B vssd1 vssd1 vccd1 vccd1 _2580_/A sky130_fd_sc_hd__and2_1
X_5298_ _5298_/A _2496_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
X_4318_ _4318_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _4326_/A sky130_fd_sc_hd__or2_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4249_ _5007_/Q _4220_/X _4247_/Y _4248_/X _4187_/X vssd1 vssd1 vccd1 vccd1 _5007_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3620_ _3590_/B _3617_/X _3619_/X vssd1 vssd1 vccd1 vccd1 _3625_/A sky130_fd_sc_hd__a21o_1
X_3551_ _3551_/A vssd1 vssd1 vccd1 vccd1 _3551_/X sky130_fd_sc_hd__clkbuf_2
X_2502_ _2503_/A vssd1 vssd1 vccd1 vccd1 _2502_/Y sky130_fd_sc_hd__inv_2
X_3482_ _4923_/Q _5091_/Q vssd1 vssd1 vccd1 vccd1 _3483_/B sky130_fd_sc_hd__and2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2433_ _2435_/A vssd1 vssd1 vccd1 vccd1 _2433_/Y sky130_fd_sc_hd__inv_2
X_5221_ _5221_/A _2421_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
X_5133__40 vssd1 vssd1 vccd1 vccd1 _5133__40/HI _5228_/A sky130_fd_sc_hd__conb_1
X_4103_ _4103_/A _4103_/B vssd1 vssd1 vccd1 vccd1 _4103_/Y sky130_fd_sc_hd__nand2_1
X_5083_ _5085_/CLK _5083_/D vssd1 vssd1 vccd1 vccd1 _5083_/Q sky130_fd_sc_hd__dfxtp_1
X_4034_ _4043_/A vssd1 vssd1 vccd1 vccd1 _4034_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _5117_/CLK _4936_/D vssd1 vssd1 vccd1 vccd1 _4936_/Q sky130_fd_sc_hd__dfxtp_1
X_4867_ _5048_/CLK _4867_/D vssd1 vssd1 vccd1 vccd1 _4867_/Q sky130_fd_sc_hd__dfxtp_1
X_3818_ _4952_/Q _3745_/X _3817_/X _3797_/X vssd1 vssd1 vccd1 vccd1 _4952_/D sky130_fd_sc_hd__o211a_1
X_4798_ _5026_/CLK _4798_/D vssd1 vssd1 vccd1 vccd1 _4798_/Q sky130_fd_sc_hd__dfxtp_1
X_3749_ _3755_/A vssd1 vssd1 vccd1 vccd1 _3749_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2982_ _2982_/A vssd1 vssd1 vccd1 vccd1 _4733_/A sky130_fd_sc_hd__buf_2
X_4721_ _4730_/A _4721_/B vssd1 vssd1 vccd1 vccd1 _4722_/A sky130_fd_sc_hd__and2_1
X_4652_ _4918_/Q _5098_/Q _4665_/S vssd1 vssd1 vccd1 vccd1 _4653_/B sky130_fd_sc_hd__mux2_1
X_3603_ _4937_/Q _5105_/Q vssd1 vssd1 vccd1 vccd1 _3603_/Y sky130_fd_sc_hd__nor2_1
X_4583_ _4592_/A _4583_/B vssd1 vssd1 vccd1 vccd1 _4584_/A sky130_fd_sc_hd__and2_1
X_3534_ _4929_/Q _5097_/Q vssd1 vssd1 vccd1 vccd1 _3535_/B sky130_fd_sc_hd__nand2_1
X_3465_ _3466_/A _3466_/B vssd1 vssd1 vccd1 vccd1 _3465_/X sky130_fd_sc_hd__or2_1
X_2416_ _2540_/A vssd1 vssd1 vccd1 vccd1 _2548_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3396_ _4910_/Q _5078_/Q _3395_/X _3388_/B vssd1 vssd1 vccd1 vccd1 _3396_/X sky130_fd_sc_hd__a31o_1
XFILLER_84_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5066_ _5066_/CLK _5066_/D vssd1 vssd1 vccd1 vccd1 _5066_/Q sky130_fd_sc_hd__dfxtp_1
X_4017_ _4017_/A vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__inv_2
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4919_ _5107_/CLK _4919_/D vssd1 vssd1 vccd1 vccd1 _4919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3250_ _3241_/A _3245_/X _3248_/X _3182_/X vssd1 vssd1 vccd1 vccd1 _3250_/X sky130_fd_sc_hd__a31o_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3181_ _3181_/A _3181_/B vssd1 vssd1 vccd1 vccd1 _3181_/Y sky130_fd_sc_hd__nand2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2965_ _3168_/B _2965_/B vssd1 vssd1 vccd1 vccd1 _2966_/B sky130_fd_sc_hd__and2_1
X_4704_ _4713_/A _4704_/B vssd1 vssd1 vccd1 vccd1 _4705_/A sky130_fd_sc_hd__and2_1
X_2896_ _2889_/X input26/X _2883_/X vssd1 vssd1 vccd1 vccd1 _2896_/X sky130_fd_sc_hd__a21bo_1
XFILLER_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4635_ _4644_/A _4635_/B vssd1 vssd1 vccd1 vccd1 _4636_/A sky130_fd_sc_hd__and2_1
X_4566_ _4575_/A _4566_/B vssd1 vssd1 vccd1 vccd1 _4567_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5117_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3517_ _3517_/A _5095_/Q vssd1 vssd1 vccd1 vccd1 _3517_/X sky130_fd_sc_hd__or2_1
XFILLER_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4497_ _4497_/A vssd1 vssd1 vccd1 vccd1 _5053_/D sky130_fd_sc_hd__clkbuf_1
X_3448_ _4906_/Q _3448_/B vssd1 vssd1 vccd1 vccd1 _3448_/X sky130_fd_sc_hd__or2_1
X_3379_ _4910_/Q _5078_/Q vssd1 vssd1 vccd1 vccd1 _3381_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5118_ _5121_/CLK _5118_/D vssd1 vssd1 vccd1 vccd1 _5118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5049_ _5062_/CLK _5049_/D vssd1 vssd1 vccd1 vccd1 _5049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2750_ _2750_/A _2750_/B vssd1 vssd1 vccd1 vccd1 _2751_/A sky130_fd_sc_hd__and2_1
X_2681_ _2681_/A vssd1 vssd1 vccd1 vccd1 _2696_/A sky130_fd_sc_hd__clkbuf_2
X_4420_ _4454_/A vssd1 vssd1 vccd1 vccd1 _4435_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4351_ _4376_/A _4351_/B vssd1 vssd1 vccd1 vccd1 _4351_/X sky130_fd_sc_hd__xor2_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ _3287_/A _3287_/B _3293_/Y _3301_/X vssd1 vssd1 vccd1 vccd1 _3303_/B sky130_fd_sc_hd__a31o_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4282_ _5011_/Q _4259_/X _4279_/Y _4280_/X _4281_/X vssd1 vssd1 vccd1 vccd1 _5011_/D
+ sky130_fd_sc_hd__o221a_1
X_3233_ _3233_/A _3233_/B _3233_/C vssd1 vssd1 vccd1 vccd1 _3233_/X sky130_fd_sc_hd__and3_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3164_ _4883_/Q _5051_/Q vssd1 vssd1 vccd1 vccd1 _3164_/X sky130_fd_sc_hd__xor2_1
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3095_ _3093_/X _3094_/Y _3078_/X vssd1 vssd1 vccd1 vccd1 _3095_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3997_ _3997_/A _3997_/B vssd1 vssd1 vccd1 vccd1 _3997_/Y sky130_fd_sc_hd__nor2_1
X_2948_ _2951_/A _2948_/B vssd1 vssd1 vccd1 vccd1 _2949_/A sky130_fd_sc_hd__and2_1
X_4618_ _4618_/A vssd1 vssd1 vccd1 vccd1 _5088_/D sky130_fd_sc_hd__clkbuf_1
X_2879_ _2862_/X input7/X _2863_/X vssd1 vssd1 vccd1 vccd1 _2879_/X sky130_fd_sc_hd__o21a_1
X_4549_ _4549_/A vssd1 vssd1 vccd1 vccd1 _5068_/D sky130_fd_sc_hd__clkbuf_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3920_ _4978_/Q _4758_/Q vssd1 vssd1 vccd1 vccd1 _3921_/B sky130_fd_sc_hd__and2_1
X_3851_ _4958_/Q vssd1 vssd1 vccd1 vccd1 _3851_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3782_ _4948_/Q _3830_/B vssd1 vssd1 vccd1 vccd1 _3782_/X sky130_fd_sc_hd__or2_1
X_2802_ _5013_/Q _4805_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _2803_/B sky130_fd_sc_hd__mux2_1
X_2733_ _2733_/A _2733_/B vssd1 vssd1 vccd1 vccd1 _2734_/A sky130_fd_sc_hd__and2_1
X_2664_ _2681_/A vssd1 vssd1 vccd1 vccd1 _2679_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4403_ _4831_/Q _4819_/Q vssd1 vssd1 vccd1 vccd1 _4403_/Y sky130_fd_sc_hd__xnor2_1
X_2595_ _4954_/Q _4746_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _2596_/B sky130_fd_sc_hd__mux2_1
X_4334_ _4335_/A _4335_/B vssd1 vssd1 vccd1 vccd1 _4336_/A sky130_fd_sc_hd__or2_1
XFILLER_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4265_ _4264_/A _4284_/B _4230_/X vssd1 vssd1 vccd1 vccd1 _4265_/X sky130_fd_sc_hd__a21o_1
X_4196_ _4196_/A _4196_/B vssd1 vssd1 vccd1 vccd1 _4198_/B sky130_fd_sc_hd__and2_1
X_3216_ _3215_/A _3233_/B _3182_/X vssd1 vssd1 vccd1 vccd1 _3216_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3147_ _3145_/X _3146_/Y _3084_/X vssd1 vssd1 vccd1 vccd1 _3147_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3078_ _3084_/A vssd1 vssd1 vccd1 vccd1 _3078_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5099_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4050_ _4051_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _4050_/X sky130_fd_sc_hd__or2_1
Xinput6 io_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_3001_ _4863_/Q _5031_/Q vssd1 vssd1 vccd1 vccd1 _3003_/A sky130_fd_sc_hd__nor2_1
X_5202__109 vssd1 vssd1 vccd1 vccd1 _5202__109/HI _5310_/A sky130_fd_sc_hd__conb_1
X_4952_ _4954_/CLK _4952_/D vssd1 vssd1 vccd1 vccd1 _4952_/Q sky130_fd_sc_hd__dfxtp_1
X_3903_ _4974_/Q _4754_/Q _3903_/C vssd1 vssd1 vccd1 vccd1 _3903_/X sky130_fd_sc_hd__and3_1
X_4883_ _5062_/CLK _4883_/D vssd1 vssd1 vccd1 vccd1 _4883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3834_ _3827_/B _3832_/Y _3833_/Y vssd1 vssd1 vccd1 vccd1 _3834_/X sky130_fd_sc_hd__o21a_1
X_3765_ _3765_/A _3765_/B vssd1 vssd1 vccd1 vccd1 _3765_/Y sky130_fd_sc_hd__nand2_1
X_2716_ _2716_/A vssd1 vssd1 vccd1 vccd1 _4780_/D sky130_fd_sc_hd__clkbuf_1
X_3696_ _3692_/Y _3712_/B _3651_/A vssd1 vssd1 vccd1 vccd1 _3696_/Y sky130_fd_sc_hd__o21ai_1
X_2647_ _2681_/A vssd1 vssd1 vccd1 vccd1 _2662_/A sky130_fd_sc_hd__clkbuf_2
X_2578_ _4949_/Q _4741_/Q _2587_/S vssd1 vssd1 vccd1 vccd1 _2579_/B sky130_fd_sc_hd__mux2_1
X_5297_ _5297_/A _2495_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
X_4317_ _4820_/Q _4808_/Q vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4248_ _4239_/A _4241_/Y _4246_/Y _4230_/X vssd1 vssd1 vccd1 vccd1 _4248_/X sky130_fd_sc_hd__a31o_1
X_4179_ _4190_/A _4161_/B _4169_/A _4189_/A _4178_/Y vssd1 vssd1 vccd1 vccd1 _4179_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3550_ _3541_/B _3547_/X _3548_/X _3467_/A vssd1 vssd1 vccd1 vccd1 _3550_/X sky130_fd_sc_hd__a31o_1
X_2501_ _2503_/A vssd1 vssd1 vccd1 vccd1 _2501_/Y sky130_fd_sc_hd__inv_2
X_5220_ _5220_/A _2420_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
X_3481_ _4923_/Q _5091_/Q vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__nor2_1
X_2432_ _2435_/A vssd1 vssd1 vccd1 vccd1 _2432_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4102_ _4103_/A _4103_/B vssd1 vssd1 vccd1 vccd1 _4102_/X sky130_fd_sc_hd__or2_1
X_5082_ _5085_/CLK _5082_/D vssd1 vssd1 vccd1 vccd1 _5082_/Q sky130_fd_sc_hd__dfxtp_1
X_4033_ _4117_/B vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4935_ _5117_/CLK _4935_/D vssd1 vssd1 vccd1 vccd1 _4935_/Q sky130_fd_sc_hd__dfxtp_1
X_4866_ _5046_/CLK _4866_/D vssd1 vssd1 vccd1 vccd1 _4866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4797_ _5004_/CLK _4797_/D vssd1 vssd1 vccd1 vccd1 _4797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3817_ _3815_/X _3816_/Y _3755_/X vssd1 vssd1 vccd1 vccd1 _3817_/X sky130_fd_sc_hd__a21o_1
X_3748_ _4129_/A _3936_/B vssd1 vssd1 vccd1 vccd1 _3755_/A sky130_fd_sc_hd__or2_2
X_3679_ _3671_/A _3673_/Y _3678_/Y vssd1 vssd1 vccd1 vccd1 _3679_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2981_ _2977_/X _2987_/A _2980_/X vssd1 vssd1 vccd1 vccd1 _2981_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4720_ _4938_/Q _5118_/Q _4732_/S vssd1 vssd1 vccd1 vccd1 _4721_/B sky130_fd_sc_hd__mux2_1
X_4651_ _4702_/A vssd1 vssd1 vccd1 vccd1 _4665_/S sky130_fd_sc_hd__clkbuf_4
Xinput20 la1_data_in[22] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_2
X_3602_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3602_/Y sky130_fd_sc_hd__inv_2
X_4582_ _4898_/Q _5078_/Q _4595_/S vssd1 vssd1 vccd1 vccd1 _4583_/B sky130_fd_sc_hd__mux2_1
X_3533_ _4929_/Q _5097_/Q vssd1 vssd1 vccd1 vccd1 _3533_/Y sky130_fd_sc_hd__nor2_1
X_3464_ _4921_/Q _5089_/Q vssd1 vssd1 vccd1 vccd1 _3466_/B sky130_fd_sc_hd__xnor2_1
X_2415_ input1/X vssd1 vssd1 vccd1 vccd1 _2540_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5208__115 vssd1 vssd1 vccd1 vccd1 _5208__115/HI _5316_/A sky130_fd_sc_hd__conb_1
X_3395_ _4911_/Q _5079_/Q vssd1 vssd1 vccd1 vccd1 _3395_/X sky130_fd_sc_hd__or2_1
XFILLER_69_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5065_ _5066_/CLK _5065_/D vssd1 vssd1 vccd1 vccd1 _5065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4016_ _4016_/A _4016_/B vssd1 vssd1 vccd1 vccd1 _4017_/A sky130_fd_sc_hd__and2_1
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4918_ _5098_/CLK _4918_/D vssd1 vssd1 vccd1 vccd1 _4918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4849_ _5041_/CLK _4849_/D vssd1 vssd1 vccd1 vccd1 _4849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _3181_/A _3181_/B vssd1 vssd1 vccd1 vccd1 _3180_/X sky130_fd_sc_hd__or2_1
XFILLER_66_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2964_ _2964_/A vssd1 vssd1 vccd1 vccd1 _4845_/D sky130_fd_sc_hd__clkbuf_1
X_4703_ _4933_/Q _5113_/Q _4716_/S vssd1 vssd1 vccd1 vccd1 _4704_/B sky130_fd_sc_hd__mux2_1
X_2895_ _2886_/X input11/X _2887_/X vssd1 vssd1 vccd1 vccd1 _2895_/X sky130_fd_sc_hd__o21a_1
X_4634_ _4913_/Q _5093_/Q _4648_/S vssd1 vssd1 vccd1 vccd1 _4635_/B sky130_fd_sc_hd__mux2_1
X_4565_ _4893_/Q _5073_/Q _4578_/S vssd1 vssd1 vccd1 vccd1 _4566_/B sky130_fd_sc_hd__mux2_1
X_3516_ _3517_/A _5095_/Q vssd1 vssd1 vccd1 vccd1 _3516_/Y sky130_fd_sc_hd__nand2_1
X_4496_ _4505_/A _4496_/B vssd1 vssd1 vccd1 vccd1 _4497_/A sky130_fd_sc_hd__and2_1
X_3447_ _3447_/A _3447_/B vssd1 vssd1 vccd1 vccd1 _3447_/X sky130_fd_sc_hd__xor2_1
X_3378_ _3372_/A _3372_/B _3377_/Y vssd1 vssd1 vccd1 vccd1 _3383_/A sky130_fd_sc_hd__o21ai_1
XFILLER_84_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5117_ _5117_/CLK _5117_/D vssd1 vssd1 vccd1 vccd1 _5117_/Q sky130_fd_sc_hd__dfxtp_1
X_5048_ _5048_/CLK _5048_/D vssd1 vssd1 vccd1 vccd1 _5048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5184__91 vssd1 vssd1 vccd1 vccd1 _5184__91/HI _5292_/A sky130_fd_sc_hd__conb_1
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2680_ _2680_/A vssd1 vssd1 vccd1 vccd1 _4770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _4335_/A _4335_/B _4341_/Y _4349_/X vssd1 vssd1 vccd1 vccd1 _4351_/B sky130_fd_sc_hd__a31o_1
X_3301_ _4898_/Q _5066_/Q _3300_/X _3293_/B vssd1 vssd1 vccd1 vccd1 _3301_/X sky130_fd_sc_hd__a31o_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4281_ _4281_/A vssd1 vssd1 vccd1 vccd1 _4281_/X sky130_fd_sc_hd__buf_2
X_3232_ _3232_/A _3232_/B _3232_/C _3236_/C vssd1 vssd1 vccd1 vccd1 _3233_/C sky130_fd_sc_hd__and4_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _3144_/A _3146_/Y _3152_/B _3160_/A _3150_/Y vssd1 vssd1 vccd1 vccd1 _3163_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3094_ _3094_/A _3094_/B vssd1 vssd1 vccd1 vccd1 _3094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3996_ _3996_/A _3996_/B _3996_/C vssd1 vssd1 vccd1 vccd1 _3997_/B sky130_fd_sc_hd__or3_1
X_2947_ _5282_/A _4857_/Q _2954_/S vssd1 vssd1 vccd1 vccd1 _2948_/B sky130_fd_sc_hd__mux2_1
X_4617_ _4626_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _4618_/A sky130_fd_sc_hd__and2_1
X_2878_ _2878_/A vssd1 vssd1 vccd1 vccd1 _2878_/X sky130_fd_sc_hd__clkbuf_2
X_4548_ _4557_/A _4548_/B vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__and2_1
XFILLER_1_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4479_ _4488_/A _4479_/B vssd1 vssd1 vccd1 vccd1 _4480_/A sky130_fd_sc_hd__and2_1
XFILLER_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3850_ _4957_/Q _3838_/X _3849_/X _3797_/X vssd1 vssd1 vccd1 vccd1 _4957_/D sky130_fd_sc_hd__o211a_1
X_2801_ _2801_/A vssd1 vssd1 vccd1 vccd1 _2815_/S sky130_fd_sc_hd__clkbuf_4
X_3781_ _3806_/A _3781_/B vssd1 vssd1 vccd1 vccd1 _3781_/X sky130_fd_sc_hd__xor2_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2732_ _4993_/Q _4785_/Q _2745_/S vssd1 vssd1 vccd1 vccd1 _2733_/B sky130_fd_sc_hd__mux2_1
X_2663_ _2663_/A vssd1 vssd1 vccd1 vccd1 _4765_/D sky130_fd_sc_hd__clkbuf_1
X_4402_ _4384_/A _4386_/Y _4391_/B _4399_/A _4389_/Y vssd1 vssd1 vccd1 vccd1 _4402_/Y
+ sky130_fd_sc_hd__a311oi_2
X_2594_ _4281_/A vssd1 vssd1 vccd1 vccd1 _2609_/A sky130_fd_sc_hd__buf_2
XFILLER_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4333_ _4333_/A _4333_/B vssd1 vssd1 vccd1 vccd1 _4335_/B sky130_fd_sc_hd__and2_1
XFILLER_5_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4264_ _4264_/A _4284_/B vssd1 vssd1 vccd1 vccd1 _4264_/Y sky130_fd_sc_hd__nor2_1
X_3215_ _3215_/A _3233_/B vssd1 vssd1 vccd1 vccd1 _3215_/Y sky130_fd_sc_hd__nor2_1
X_4195_ _5012_/Q _4792_/Q vssd1 vssd1 vccd1 vccd1 _4196_/B sky130_fd_sc_hd__or2_1
X_3146_ _3146_/A _3146_/B vssd1 vssd1 vccd1 vccd1 _3146_/Y sky130_fd_sc_hd__nand2_1
X_3077_ _4223_/A _3077_/B vssd1 vssd1 vccd1 vccd1 _3084_/A sky130_fd_sc_hd__or2_2
XFILLER_54_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3979_ _4973_/Q _4021_/B vssd1 vssd1 vccd1 vccd1 _3979_/X sky130_fd_sc_hd__or2_1
XFILLER_40_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5154__61 vssd1 vssd1 vccd1 vccd1 _5154__61/HI _5249_/A sky130_fd_sc_hd__conb_1
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 io_in[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3000_ _2991_/Y _2980_/X _2999_/Y _2967_/A vssd1 vssd1 vccd1 vccd1 _4850_/D sky130_fd_sc_hd__a211oi_1
XFILLER_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4951_ _4954_/CLK _4951_/D vssd1 vssd1 vccd1 vccd1 _4951_/Q sky130_fd_sc_hd__dfxtp_1
X_3902_ _3902_/A _3902_/B _3902_/C vssd1 vssd1 vccd1 vccd1 _3902_/X sky130_fd_sc_hd__and3_1
X_4882_ _5062_/CLK _4882_/D vssd1 vssd1 vccd1 vccd1 _4882_/Q sky130_fd_sc_hd__dfxtp_1
X_3833_ _4967_/Q _4747_/Q vssd1 vssd1 vccd1 vccd1 _3833_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3764_ _3765_/A _3765_/B vssd1 vssd1 vccd1 vccd1 _3764_/X sky130_fd_sc_hd__or2_1
X_2715_ _2715_/A _2715_/B vssd1 vssd1 vccd1 vccd1 _2716_/A sky130_fd_sc_hd__and2_1
X_3695_ _3693_/Y _3695_/B vssd1 vssd1 vccd1 vccd1 _3712_/B sky130_fd_sc_hd__and2b_1
X_2646_ _2646_/A vssd1 vssd1 vccd1 vccd1 _4760_/D sky130_fd_sc_hd__clkbuf_1
X_2577_ _4281_/A vssd1 vssd1 vccd1 vccd1 _2592_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5296_ _5296_/A _2494_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
X_4316_ _4820_/Q _4808_/Q vssd1 vssd1 vccd1 vccd1 _4316_/X sky130_fd_sc_hd__or2_1
XFILLER_19_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4247_ _4239_/A _4241_/Y _4246_/Y vssd1 vssd1 vccd1 vccd1 _4247_/Y sky130_fd_sc_hd__a21oi_1
X_4178_ _4177_/Y _4169_/B _4175_/Y vssd1 vssd1 vccd1 vccd1 _4178_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3129_ _4879_/Q _5047_/Q vssd1 vssd1 vccd1 vccd1 _3137_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2500_ _2503_/A vssd1 vssd1 vccd1 vccd1 _2500_/Y sky130_fd_sc_hd__inv_2
X_3480_ _3470_/Y _3461_/X _3478_/Y _3479_/X vssd1 vssd1 vccd1 vccd1 _4910_/D sky130_fd_sc_hd__a211oi_1
X_2431_ _2435_/A vssd1 vssd1 vccd1 vccd1 _2431_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4101_ _4101_/A _4101_/B vssd1 vssd1 vccd1 vccd1 _4103_/B sky130_fd_sc_hd__and2_1
X_5081_ _5091_/CLK _5081_/D vssd1 vssd1 vccd1 vccd1 _5081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4032_ _4032_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _4117_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4934_ _5114_/CLK _4934_/D vssd1 vssd1 vccd1 vccd1 _4934_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4972_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4865_ _5046_/CLK _4865_/D vssd1 vssd1 vccd1 vccd1 _4865_/Q sky130_fd_sc_hd__dfxtp_1
X_4796_ _5004_/CLK _4796_/D vssd1 vssd1 vccd1 vccd1 _4796_/Q sky130_fd_sc_hd__dfxtp_1
X_3816_ _3816_/A _3816_/B vssd1 vssd1 vccd1 vccd1 _3816_/Y sky130_fd_sc_hd__nand2_2
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3747_ _4956_/Q _4736_/Q vssd1 vssd1 vccd1 vccd1 _3754_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3678_ _3678_/A _3678_/B vssd1 vssd1 vccd1 vccd1 _3678_/Y sky130_fd_sc_hd__nor2_1
X_2629_ _2681_/A vssd1 vssd1 vccd1 vccd1 _2645_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5124__31 vssd1 vssd1 vccd1 vccd1 _5124__31/HI _5219_/A sky130_fd_sc_hd__conb_1
X_5279_ _5279_/A _2474_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2980_ _2988_/A vssd1 vssd1 vccd1 vccd1 _2980_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4650_ _4650_/A vssd1 vssd1 vccd1 vccd1 _5097_/D sky130_fd_sc_hd__clkbuf_1
Xinput10 io_in[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_2
Xinput21 la1_data_in[23] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_2
X_3601_ _4938_/Q _5106_/Q vssd1 vssd1 vccd1 vccd1 _3616_/A sky130_fd_sc_hd__xor2_2
X_4581_ _4615_/A vssd1 vssd1 vccd1 vccd1 _4595_/S sky130_fd_sc_hd__clkbuf_2
X_3532_ _4916_/Q _3457_/X _3531_/X _3503_/X vssd1 vssd1 vccd1 vccd1 _4916_/D sky130_fd_sc_hd__o211a_1
XFILLER_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3463_ _4908_/Q _3457_/X _3462_/X _3434_/X vssd1 vssd1 vccd1 vccd1 _4908_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3394_ _3394_/A _3394_/B vssd1 vssd1 vccd1 vccd1 _3422_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _5070_/CLK _5064_/D vssd1 vssd1 vccd1 vccd1 _5064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4015_ _4990_/Q _4770_/Q vssd1 vssd1 vccd1 vccd1 _4016_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4917_ _5107_/CLK _4917_/D vssd1 vssd1 vccd1 vccd1 _4917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4848_ _5041_/CLK _4848_/D vssd1 vssd1 vccd1 vccd1 _4848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4779_ _4995_/CLK _4779_/D vssd1 vssd1 vccd1 vccd1 _4779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2963_ _3037_/A _4032_/A _2963_/C vssd1 vssd1 vccd1 vccd1 _2964_/A sky130_fd_sc_hd__and3_1
X_4702_ _4702_/A vssd1 vssd1 vccd1 vccd1 _4716_/S sky130_fd_sc_hd__buf_2
X_2894_ _2878_/X _4827_/Q _2892_/X _2893_/X _2876_/X vssd1 vssd1 vccd1 vccd1 _4827_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633_ _4702_/A vssd1 vssd1 vccd1 vccd1 _4648_/S sky130_fd_sc_hd__buf_2
X_4564_ _4615_/A vssd1 vssd1 vccd1 vccd1 _4578_/S sky130_fd_sc_hd__buf_2
X_3515_ _3520_/A _3507_/X _3521_/B _3521_/C vssd1 vssd1 vccd1 vccd1 _3515_/X sky130_fd_sc_hd__o2bb2a_1
X_4495_ _4873_/Q _5053_/Q _4508_/S vssd1 vssd1 vccd1 vccd1 _4496_/B sky130_fd_sc_hd__mux2_1
X_3446_ _3430_/A _3432_/Y _3438_/B _3436_/Y vssd1 vssd1 vccd1 vccd1 _3447_/B sky130_fd_sc_hd__a31o_1
X_3377_ _4909_/Q _5077_/Q vssd1 vssd1 vccd1 vccd1 _3377_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5116_ _5117_/CLK _5116_/D vssd1 vssd1 vccd1 vccd1 _5116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5047_ _5048_/CLK _5047_/D vssd1 vssd1 vccd1 vccd1 _5047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5079_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3300_ _4899_/Q _5067_/Q vssd1 vssd1 vccd1 vccd1 _3300_/X sky130_fd_sc_hd__or2_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4280_ _4276_/Y _4270_/X _4283_/B _4285_/C _4230_/A vssd1 vssd1 vccd1 vccd1 _4280_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _4879_/Q _3223_/A _3228_/Y _3229_/X _3230_/X vssd1 vssd1 vccd1 vccd1 _4879_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _3078_/X _3160_/X _3161_/X _3148_/X vssd1 vssd1 vccd1 vccd1 _4870_/D sky130_fd_sc_hd__o211a_1
X_3093_ _3094_/A _3094_/B vssd1 vssd1 vccd1 vccd1 _3093_/X sky130_fd_sc_hd__or2_1
X_3995_ _3995_/A _3996_/C vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__or2_1
XFILLER_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2946_ _2946_/A vssd1 vssd1 vccd1 vccd1 _4840_/D sky130_fd_sc_hd__clkbuf_1
X_2877_ _2855_/X _4823_/Q _2874_/X _2875_/X _2876_/X vssd1 vssd1 vccd1 vccd1 _4823_/D
+ sky130_fd_sc_hd__o221a_1
X_4616_ _4908_/Q _5088_/Q _4629_/S vssd1 vssd1 vccd1 vccd1 _4617_/B sky130_fd_sc_hd__mux2_1
X_4547_ _4888_/Q _5068_/Q _4561_/S vssd1 vssd1 vccd1 vccd1 _4548_/B sky130_fd_sc_hd__mux2_1
X_4478_ _4868_/Q _5048_/Q _4491_/S vssd1 vssd1 vccd1 vccd1 _4479_/B sky130_fd_sc_hd__mux2_1
X_3429_ _4916_/Q _5084_/Q vssd1 vssd1 vccd1 vccd1 _3430_/B sky130_fd_sc_hd__or2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2800_ _2800_/A vssd1 vssd1 vccd1 vccd1 _4804_/D sky130_fd_sc_hd__clkbuf_1
X_3780_ _3765_/A _3765_/B _3770_/Y _3779_/X vssd1 vssd1 vccd1 vccd1 _3781_/B sky130_fd_sc_hd__a31o_1
X_2731_ _2801_/A vssd1 vssd1 vccd1 vccd1 _2745_/S sky130_fd_sc_hd__buf_2
X_2662_ _2662_/A _2662_/B vssd1 vssd1 vccd1 vccd1 _2663_/A sky130_fd_sc_hd__and2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4401_ _4319_/X _4399_/X _4400_/X _2869_/X vssd1 vssd1 vccd1 vccd1 _5026_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2593_ _2593_/A vssd1 vssd1 vccd1 vccd1 _4745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4332_ _4822_/Q _4810_/Q vssd1 vssd1 vccd1 vccd1 _4333_/B sky130_fd_sc_hd__or2_1
X_4263_ _4263_/A _4263_/B vssd1 vssd1 vccd1 vccd1 _4284_/B sky130_fd_sc_hd__and2_1
X_3214_ _3212_/Y _3214_/B vssd1 vssd1 vccd1 vccd1 _3233_/B sky130_fd_sc_hd__and2b_1
X_4194_ _5012_/Q _4792_/Q vssd1 vssd1 vccd1 vccd1 _4196_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3145_ _3146_/A _3146_/B vssd1 vssd1 vccd1 vccd1 _3145_/X sky130_fd_sc_hd__or2_1
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3076_ _4872_/Q _5040_/Q vssd1 vssd1 vccd1 vccd1 _3083_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ _3978_/A _3997_/A vssd1 vssd1 vccd1 vccd1 _3978_/X sky130_fd_sc_hd__xor2_1
X_2929_ _2954_/S vssd1 vssd1 vccd1 vccd1 _2944_/S sky130_fd_sc_hd__buf_2
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 io_in[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4950_ _4954_/CLK _4950_/D vssd1 vssd1 vccd1 vccd1 _4950_/Q sky130_fd_sc_hd__dfxtp_1
X_3901_ _3901_/A _3901_/B _3903_/C vssd1 vssd1 vccd1 vccd1 _3902_/C sky130_fd_sc_hd__and3_1
X_4881_ _5099_/CLK _4881_/D vssd1 vssd1 vccd1 vccd1 _4881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3832_ _3814_/A _3816_/Y _3821_/B _3829_/A _3819_/Y vssd1 vssd1 vccd1 vccd1 _3832_/Y
+ sky130_fd_sc_hd__a311oi_2
X_3763_ _3763_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3765_/B sky130_fd_sc_hd__and2_1
X_2714_ _4988_/Q _4780_/Q _2727_/S vssd1 vssd1 vccd1 vccd1 _2715_/B sky130_fd_sc_hd__mux2_1
X_3694_ _5117_/Q _4949_/Q vssd1 vssd1 vccd1 vccd1 _3695_/B sky130_fd_sc_hd__nand2_1
X_2645_ _2645_/A _2645_/B vssd1 vssd1 vccd1 vccd1 _2646_/A sky130_fd_sc_hd__and2_1
XFILLER_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2576_ _2576_/A vssd1 vssd1 vccd1 vccd1 _4740_/D sky130_fd_sc_hd__clkbuf_1
X_4315_ _4400_/B vssd1 vssd1 vccd1 vccd1 _4315_/X sky130_fd_sc_hd__clkbuf_2
X_5295_ _5295_/A _2493_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
X_4246_ _4246_/A _4246_/B vssd1 vssd1 vccd1 vccd1 _4246_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4177_ _5008_/Q _4788_/Q vssd1 vssd1 vccd1 vccd1 _4177_/Y sky130_fd_sc_hd__nand2_1
X_3128_ _4878_/Q _5046_/Q vssd1 vssd1 vccd1 vccd1 _3128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3059_ _3059_/A _3059_/B vssd1 vssd1 vccd1 vccd1 _3061_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2430_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2435_/A sky130_fd_sc_hd__buf_12
X_4100_ _5000_/Q _4780_/Q vssd1 vssd1 vccd1 vccd1 _4101_/B sky130_fd_sc_hd__or2_1
X_5080_ _5091_/CLK _5080_/D vssd1 vssd1 vccd1 vccd1 _5080_/Q sky130_fd_sc_hd__dfxtp_1
X_4031_ _4223_/B vssd1 vssd1 vccd1 vccd1 _4318_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4933_ _5117_/CLK _4933_/D vssd1 vssd1 vccd1 vccd1 _4933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4864_ _5048_/CLK _4864_/D vssd1 vssd1 vccd1 vccd1 _4864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4795_ _5010_/CLK _4795_/D vssd1 vssd1 vccd1 vccd1 _4795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3815_ _3816_/A _3816_/B vssd1 vssd1 vccd1 vccd1 _3815_/X sky130_fd_sc_hd__or2_1
X_3746_ _4956_/Q _4736_/Q vssd1 vssd1 vccd1 vccd1 _3746_/X sky130_fd_sc_hd__or2_1
X_3677_ _5115_/Q _4947_/Q vssd1 vssd1 vccd1 vccd1 _3678_/B sky130_fd_sc_hd__and2_1
X_2628_ _2628_/A vssd1 vssd1 vccd1 vccd1 _4755_/D sky130_fd_sc_hd__clkbuf_1
X_2559_ _3133_/A vssd1 vssd1 vccd1 vccd1 _4281_/A sky130_fd_sc_hd__buf_2
X_5278_ _5278_/A _2472_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
X_4229_ _4229_/A _4229_/B vssd1 vssd1 vccd1 vccd1 _4229_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput22 la1_data_in[24] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
X_4580_ _4580_/A vssd1 vssd1 vccd1 vccd1 _5077_/D sky130_fd_sc_hd__clkbuf_1
Xinput11 io_in[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_4
X_3600_ _4925_/Q _3593_/X _3598_/Y _3599_/X _3551_/X vssd1 vssd1 vccd1 vccd1 _4925_/D
+ sky130_fd_sc_hd__o221a_1
X_3531_ _3529_/Y _3530_/X _3467_/X vssd1 vssd1 vccd1 vccd1 _3531_/X sky130_fd_sc_hd__a21o_1
X_3462_ _3458_/X _3466_/A _3461_/X vssd1 vssd1 vccd1 vccd1 _3462_/X sky130_fd_sc_hd__a21o_1
X_3393_ _4912_/Q _5080_/Q vssd1 vssd1 vccd1 vccd1 _3394_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5063_ _5099_/CLK _5063_/D vssd1 vssd1 vccd1 vccd1 _5063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4014_ _4990_/Q _4770_/Q vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__or2_1
X_4916_ _5094_/CLK _4916_/D vssd1 vssd1 vccd1 vccd1 _4916_/Q sky130_fd_sc_hd__dfxtp_1
X_4847_ _5051_/CLK _4847_/D vssd1 vssd1 vccd1 vccd1 _4847_/Q sky130_fd_sc_hd__dfxtp_1
X_4778_ _4995_/CLK _4778_/D vssd1 vssd1 vccd1 vccd1 _4778_/Q sky130_fd_sc_hd__dfxtp_1
X_3729_ _3720_/A _3722_/Y _3728_/X vssd1 vssd1 vccd1 vccd1 _3729_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5026_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2962_ _3168_/B _2965_/B vssd1 vssd1 vccd1 vccd1 _2963_/C sky130_fd_sc_hd__or2_1
XFILLER_15_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4701_ _4701_/A vssd1 vssd1 vccd1 vccd1 _5112_/D sky130_fd_sc_hd__clkbuf_1
X_4632_ _4632_/A vssd1 vssd1 vccd1 vccd1 _4702_/A sky130_fd_sc_hd__clkbuf_2
X_2893_ _2889_/X input25/X _2883_/X vssd1 vssd1 vccd1 vccd1 _2893_/X sky130_fd_sc_hd__a21bo_1
X_5214__121 vssd1 vssd1 vccd1 vccd1 _5214__121/HI _5322_/A sky130_fd_sc_hd__conb_1
XFILLER_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4563_ _4563_/A vssd1 vssd1 vccd1 vccd1 _5072_/D sky130_fd_sc_hd__clkbuf_1
X_4494_ _4528_/A vssd1 vssd1 vccd1 vccd1 _4508_/S sky130_fd_sc_hd__buf_2
X_3514_ _3517_/A _5095_/Q vssd1 vssd1 vccd1 vccd1 _3521_/C sky130_fd_sc_hd__nor2_1
X_3445_ _3445_/A _3445_/B vssd1 vssd1 vccd1 vccd1 _3447_/A sky130_fd_sc_hd__or2_1
X_3376_ _4898_/Q vssd1 vssd1 vccd1 vccd1 _3376_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5115_ _5117_/CLK _5115_/D vssd1 vssd1 vccd1 vccd1 _5115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5046_ _5046_/CLK _5046_/D vssd1 vssd1 vccd1 vccd1 _5046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5175__82 vssd1 vssd1 vccd1 vccd1 _5175__82/HI _5270_/A sky130_fd_sc_hd__conb_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3551_/A vssd1 vssd1 vccd1 vccd1 _3230_/X sky130_fd_sc_hd__buf_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _4870_/Q _3161_/B vssd1 vssd1 vccd1 vccd1 _3161_/X sky130_fd_sc_hd__or2_1
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3092_ _3092_/A _3092_/B vssd1 vssd1 vccd1 vccd1 _3094_/B sky130_fd_sc_hd__and2_1
XFILLER_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3994_ _4975_/Q _3933_/A _3990_/X _3993_/X _3962_/X vssd1 vssd1 vccd1 vccd1 _4975_/D
+ sky130_fd_sc_hd__o221a_1
X_2945_ _2951_/A _2945_/B vssd1 vssd1 vccd1 vccd1 _2946_/A sky130_fd_sc_hd__and2_1
X_2876_ _3037_/A vssd1 vssd1 vccd1 vccd1 _2876_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4615_ _4615_/A vssd1 vssd1 vccd1 vccd1 _4629_/S sky130_fd_sc_hd__clkbuf_2
X_4546_ _4615_/A vssd1 vssd1 vccd1 vccd1 _4561_/S sky130_fd_sc_hd__buf_2
X_4477_ _4528_/A vssd1 vssd1 vccd1 vccd1 _4491_/S sky130_fd_sc_hd__buf_2
X_3428_ _4916_/Q _5084_/Q vssd1 vssd1 vccd1 vccd1 _3430_/A sky130_fd_sc_hd__nand2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _3349_/B _3356_/X _3357_/X _3288_/X vssd1 vssd1 vccd1 vccd1 _3359_/Y sky130_fd_sc_hd__a31oi_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5029_ _5030_/CLK _5029_/D vssd1 vssd1 vccd1 vccd1 _5029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2730_ _4719_/A vssd1 vssd1 vccd1 vccd1 _2801_/A sky130_fd_sc_hd__clkbuf_2
X_2661_ _4973_/Q _4765_/Q _2674_/S vssd1 vssd1 vccd1 vccd1 _2662_/B sky130_fd_sc_hd__mux2_1
X_4400_ _5026_/Q _4400_/B vssd1 vssd1 vccd1 vccd1 _4400_/X sky130_fd_sc_hd__or2_1
X_2592_ _2592_/A _2592_/B vssd1 vssd1 vccd1 vccd1 _2593_/A sky130_fd_sc_hd__and2_1
X_4331_ _4822_/Q _4810_/Q vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__nand2_1
X_4262_ _5021_/Q _4801_/Q vssd1 vssd1 vccd1 vccd1 _4263_/B sky130_fd_sc_hd__nand2_1
X_3213_ _4889_/Q _5057_/Q vssd1 vssd1 vccd1 vccd1 _3214_/B sky130_fd_sc_hd__nand2_1
X_4193_ _4161_/B _4190_/X _4192_/X vssd1 vssd1 vccd1 vccd1 _4198_/A sky130_fd_sc_hd__a21o_1
X_3144_ _3144_/A _3144_/B vssd1 vssd1 vccd1 vccd1 _3146_/B sky130_fd_sc_hd__and2_1
X_3075_ _4872_/Q _5040_/Q vssd1 vssd1 vccd1 vccd1 _3075_/X sky130_fd_sc_hd__or2_1
XFILLER_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3977_ _3977_/A _3976_/Y vssd1 vssd1 vccd1 vccd1 _3997_/A sky130_fd_sc_hd__or2b_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2928_ _2928_/A vssd1 vssd1 vccd1 vccd1 _4835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2859_ input2/X input3/X _2905_/A vssd1 vssd1 vccd1 vccd1 _2859_/X sky130_fd_sc_hd__or3b_1
XFILLER_2_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4529_ _4883_/Q _5063_/Q _4542_/S vssd1 vssd1 vccd1 vccd1 _4530_/B sky130_fd_sc_hd__mux2_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5145__52 vssd1 vssd1 vccd1 vccd1 _5145__52/HI _5240_/A sky130_fd_sc_hd__conb_1
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 io_in[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3900_ _4963_/Q _3878_/X _3898_/Y _3899_/X _3866_/X vssd1 vssd1 vccd1 vccd1 _4963_/D
+ sky130_fd_sc_hd__o221a_1
X_4880_ _5062_/CLK _4880_/D vssd1 vssd1 vccd1 vccd1 _4880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3831_ _3749_/X _3829_/X _3830_/X _3797_/X vssd1 vssd1 vccd1 vccd1 _4954_/D sky130_fd_sc_hd__o211a_1
X_3762_ _4958_/Q _4738_/Q vssd1 vssd1 vccd1 vccd1 _3763_/B sky130_fd_sc_hd__or2_1
X_2713_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2727_/S sky130_fd_sc_hd__clkbuf_2
X_3693_ _5117_/Q _4949_/Q vssd1 vssd1 vccd1 vccd1 _3693_/Y sky130_fd_sc_hd__nor2_1
X_2644_ _4968_/Q _4760_/Q _2657_/S vssd1 vssd1 vccd1 vccd1 _2645_/B sky130_fd_sc_hd__mux2_1
X_2575_ _2575_/A _2575_/B vssd1 vssd1 vccd1 vccd1 _2576_/A sky130_fd_sc_hd__and2_1
X_4314_ _4361_/A vssd1 vssd1 vccd1 vccd1 _4400_/B sky130_fd_sc_hd__clkbuf_1
X_5294_ _5294_/A _2490_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
X_4245_ _5019_/Q _4799_/Q vssd1 vssd1 vccd1 vccd1 _4246_/B sky130_fd_sc_hd__and2_1
X_4176_ _4170_/A _4169_/B _4174_/Y _4175_/Y vssd1 vssd1 vccd1 vccd1 _4176_/X sky130_fd_sc_hd__a211o_1
X_3127_ _4866_/Q _3074_/X _3126_/X _3063_/X vssd1 vssd1 vccd1 vccd1 _4866_/D sky130_fd_sc_hd__o211a_1
XFILLER_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3058_ _4870_/Q _5038_/Q vssd1 vssd1 vccd1 vccd1 _3059_/B sky130_fd_sc_hd__nand2_1
XFILLER_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4030_ _4847_/Q _4030_/B vssd1 vssd1 vccd1 vccd1 _4223_/B sky130_fd_sc_hd__or2_1
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4932_ _5117_/CLK _4932_/D vssd1 vssd1 vccd1 vccd1 _4932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4863_ _5046_/CLK _4863_/D vssd1 vssd1 vccd1 vccd1 _4863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4794_ _5010_/CLK _4794_/D vssd1 vssd1 vccd1 vccd1 _4794_/Q sky130_fd_sc_hd__dfxtp_1
X_3814_ _3814_/A _3814_/B vssd1 vssd1 vccd1 vccd1 _3816_/B sky130_fd_sc_hd__and2_1
XFILLER_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3745_ _3830_/B vssd1 vssd1 vccd1 vccd1 _3745_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3676_ _5115_/Q _4947_/Q vssd1 vssd1 vccd1 vccd1 _3678_/A sky130_fd_sc_hd__nor2_1
X_2627_ _2627_/A _2627_/B vssd1 vssd1 vccd1 vccd1 _2628_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5107_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2558_ _2558_/A vssd1 vssd1 vccd1 vccd1 _4735_/D sky130_fd_sc_hd__clkbuf_1
X_5277_ _5277_/A _2471_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
X_2489_ _2490_/A vssd1 vssd1 vccd1 vccd1 _2489_/Y sky130_fd_sc_hd__inv_2
X_4228_ _4229_/A _4229_/B vssd1 vssd1 vccd1 vccd1 _4228_/X sky130_fd_sc_hd__or2_1
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4159_ _5006_/Q _4786_/Q _4158_/X _4151_/B vssd1 vssd1 vccd1 vccd1 _4159_/X sky130_fd_sc_hd__a31o_1
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 io_in[20] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput23 la1_data_in[25] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
X_3530_ _3529_/A _3529_/B _3529_/C vssd1 vssd1 vccd1 vccd1 _3530_/X sky130_fd_sc_hd__a21o_1
X_3461_ _3467_/A vssd1 vssd1 vccd1 vccd1 _3461_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3392_ _4912_/Q _5080_/Q vssd1 vssd1 vccd1 vccd1 _3394_/A sky130_fd_sc_hd__and2_1
X_5062_ _5062_/CLK _5062_/D vssd1 vssd1 vccd1 vccd1 _5062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4013_ _4977_/Q _3933_/A _4011_/Y _4012_/X _3962_/X vssd1 vssd1 vccd1 vccd1 _4977_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_80_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4915_ _5107_/CLK _4915_/D vssd1 vssd1 vccd1 vccd1 _4915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4846_ _5051_/CLK _4846_/D vssd1 vssd1 vccd1 vccd1 _4846_/Q sky130_fd_sc_hd__dfxtp_1
X_4777_ _4995_/CLK _4777_/D vssd1 vssd1 vccd1 vccd1 _4777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3728_ _3726_/Y _3728_/B vssd1 vssd1 vccd1 vccd1 _3728_/X sky130_fd_sc_hd__and2b_1
X_3659_ _3945_/A vssd1 vssd1 vccd1 vccd1 _3659_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2961_ _4037_/A vssd1 vssd1 vccd1 vccd1 _4032_/A sky130_fd_sc_hd__buf_2
X_4700_ _4713_/A _4700_/B vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__and2_1
X_4631_ _4631_/A vssd1 vssd1 vccd1 vccd1 _5092_/D sky130_fd_sc_hd__clkbuf_1
X_2892_ _2886_/X input10/X _2887_/X vssd1 vssd1 vccd1 vccd1 _2892_/X sky130_fd_sc_hd__o21a_1
X_4562_ _4575_/A _4562_/B vssd1 vssd1 vccd1 vccd1 _4563_/A sky130_fd_sc_hd__and2_1
X_4493_ _4493_/A vssd1 vssd1 vccd1 vccd1 _5052_/D sky130_fd_sc_hd__clkbuf_1
X_3513_ _4927_/Q vssd1 vssd1 vccd1 vccd1 _3517_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3444_ _4918_/Q _5086_/Q vssd1 vssd1 vccd1 vccd1 _3445_/B sky130_fd_sc_hd__and2_1
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3375_ _4897_/Q _3363_/X _3374_/X _3353_/X vssd1 vssd1 vccd1 vccd1 _4897_/D sky130_fd_sc_hd__o211a_1
X_5114_ _5114_/CLK _5114_/D vssd1 vssd1 vccd1 vccd1 _5114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5045_ _5046_/CLK _5045_/D vssd1 vssd1 vccd1 vccd1 _5045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_43_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5048_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4829_ _4836_/CLK _4829_/D vssd1 vssd1 vccd1 vccd1 _4829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5196__103 vssd1 vssd1 vccd1 vccd1 _5196__103/HI _5304_/A sky130_fd_sc_hd__conb_1
XFILLER_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5190__97 vssd1 vssd1 vccd1 vccd1 _5190__97/HI _5298_/A sky130_fd_sc_hd__conb_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3160_/A _3160_/B vssd1 vssd1 vccd1 vccd1 _3160_/X sky130_fd_sc_hd__xor2_1
X_3091_ _4874_/Q _5042_/Q vssd1 vssd1 vccd1 vccd1 _3092_/B sky130_fd_sc_hd__or2_1
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3993_ _3995_/A _3983_/X _3991_/Y _3992_/X _3943_/A vssd1 vssd1 vccd1 vccd1 _3993_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2944_ _5281_/A _4856_/Q _2944_/S vssd1 vssd1 vccd1 vccd1 _2945_/B sky130_fd_sc_hd__mux2_1
X_2875_ _2865_/X input21/X _2878_/A vssd1 vssd1 vccd1 vccd1 _2875_/X sky130_fd_sc_hd__a21bo_1
X_4614_ _4614_/A vssd1 vssd1 vccd1 vccd1 _5087_/D sky130_fd_sc_hd__clkbuf_1
X_4545_ _4632_/A vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__clkbuf_2
X_4476_ _4476_/A vssd1 vssd1 vccd1 vccd1 _5047_/D sky130_fd_sc_hd__clkbuf_1
X_3427_ _3398_/B _3422_/X _3426_/X vssd1 vssd1 vccd1 vccd1 _3432_/A sky130_fd_sc_hd__a21o_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _3349_/B _3356_/X _3357_/X vssd1 vssd1 vccd1 vccd1 _3358_/X sky130_fd_sc_hd__a21o_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _3286_/X _3287_/Y _3288_/X vssd1 vssd1 vccd1 vccd1 _3289_/X sky130_fd_sc_hd__a21o_1
X_5028_ _5030_/CLK _5028_/D vssd1 vssd1 vccd1 vccd1 _5028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2660_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2674_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2591_ _4953_/Q _4745_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _2592_/B sky130_fd_sc_hd__mux2_1
X_4330_ _4325_/A _4325_/B _4329_/Y vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__o21ai_1
X_4261_ _5021_/Q _4801_/Q vssd1 vssd1 vccd1 vccd1 _4263_/A sky130_fd_sc_hd__or2_1
X_3212_ _4889_/Q _5057_/Q vssd1 vssd1 vccd1 vccd1 _3212_/Y sky130_fd_sc_hd__nor2_1
X_4192_ _5011_/Q _4791_/Q _4178_/Y _4190_/C _4191_/X vssd1 vssd1 vccd1 vccd1 _4192_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3143_ _4880_/Q _5048_/Q vssd1 vssd1 vccd1 vccd1 _3144_/B sky130_fd_sc_hd__or2_1
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3074_ _3074_/A vssd1 vssd1 vccd1 vccd1 _3074_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3976_ _4985_/Q _4765_/Q vssd1 vssd1 vccd1 vccd1 _3976_/Y sky130_fd_sc_hd__nand2_1
X_2927_ _2934_/A _2927_/B vssd1 vssd1 vccd1 vccd1 _2928_/A sky130_fd_sc_hd__and2_1
X_2858_ _2905_/A _2858_/B _2889_/A vssd1 vssd1 vccd1 vccd1 _2858_/X sky130_fd_sc_hd__or3b_1
X_2789_ _5009_/Q _4801_/Q _2798_/S vssd1 vssd1 vccd1 vccd1 _2790_/B sky130_fd_sc_hd__mux2_1
X_4528_ _4528_/A vssd1 vssd1 vccd1 vccd1 _4542_/S sky130_fd_sc_hd__clkbuf_4
X_4459_ _4528_/A vssd1 vssd1 vccd1 vccd1 _4474_/S sky130_fd_sc_hd__buf_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5160__67 vssd1 vssd1 vccd1 vccd1 _5160__67/HI _5255_/A sky130_fd_sc_hd__conb_1
XFILLER_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3830_ _4954_/Q _3830_/B vssd1 vssd1 vccd1 vccd1 _3830_/X sky130_fd_sc_hd__or2_1
X_3761_ _4958_/Q _4738_/Q vssd1 vssd1 vccd1 vccd1 _3763_/A sky130_fd_sc_hd__nand2_1
X_2712_ _2712_/A vssd1 vssd1 vccd1 vccd1 _4779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3692_ _3712_/A _3689_/B _3685_/A vssd1 vssd1 vccd1 vccd1 _3692_/Y sky130_fd_sc_hd__a21oi_1
X_2643_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2657_/S sky130_fd_sc_hd__buf_2
X_2574_ _4948_/Q _4740_/Q _2587_/S vssd1 vssd1 vccd1 vccd1 _2575_/B sky130_fd_sc_hd__mux2_1
X_4313_ _4318_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _4361_/A sky130_fd_sc_hd__nor2_1
X_5293_ _5293_/A _2489_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4244_ _5019_/Q _4799_/Q vssd1 vssd1 vccd1 vccd1 _4246_/A sky130_fd_sc_hd__nor2_1
X_4175_ _5009_/Q _4789_/Q vssd1 vssd1 vccd1 vccd1 _4175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3126_ _3122_/X _3125_/X _3084_/X vssd1 vssd1 vccd1 vccd1 _3126_/X sky130_fd_sc_hd__a21o_1
XFILLER_82_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3057_ _4870_/Q _5038_/Q vssd1 vssd1 vccd1 vccd1 _3059_/A sky130_fd_sc_hd__or2_1
XFILLER_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _3959_/A _3959_/B vssd1 vssd1 vccd1 vccd1 _3959_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4931_ _5121_/CLK _4931_/D vssd1 vssd1 vccd1 vccd1 _4931_/Q sky130_fd_sc_hd__dfxtp_1
X_4862_ _5046_/CLK _4862_/D vssd1 vssd1 vccd1 vccd1 _4862_/Q sky130_fd_sc_hd__dfxtp_1
X_3813_ _4964_/Q _4744_/Q vssd1 vssd1 vccd1 vccd1 _3814_/B sky130_fd_sc_hd__or2_1
X_4793_ _4999_/CLK _4793_/D vssd1 vssd1 vccd1 vccd1 _4793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3744_ _4125_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _3830_/B sky130_fd_sc_hd__nor2_2
X_3675_ _3666_/Y _3656_/X _3674_/Y _3479_/X vssd1 vssd1 vccd1 vccd1 _4934_/D sky130_fd_sc_hd__a211oi_1
X_2626_ _4963_/Q _4755_/Q _2639_/S vssd1 vssd1 vccd1 vccd1 _2627_/B sky130_fd_sc_hd__mux2_1
X_2557_ _2557_/A _2557_/B vssd1 vssd1 vccd1 vccd1 _2558_/A sky130_fd_sc_hd__and2_1
X_5276_ _5276_/A _2470_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
X_2488_ _2490_/A vssd1 vssd1 vccd1 vccd1 _2488_/Y sky130_fd_sc_hd__inv_2
X_4227_ _5017_/Q _4797_/Q vssd1 vssd1 vccd1 vccd1 _4229_/B sky130_fd_sc_hd__xnor2_1
XFILLER_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4158_ _5007_/Q _4787_/Q vssd1 vssd1 vccd1 vccd1 _4158_/X sky130_fd_sc_hd__or2_1
XFILLER_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4089_ _4084_/Y _4086_/X _4092_/B _4096_/C vssd1 vssd1 vccd1 vccd1 _4089_/Y sky130_fd_sc_hd__a22oi_1
X_3109_ _3138_/A _3109_/B vssd1 vssd1 vccd1 vccd1 _3109_/X sky130_fd_sc_hd__xor2_1
XFILLER_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130__37 vssd1 vssd1 vccd1 vccd1 _5130__37/HI _5225_/A sky130_fd_sc_hd__conb_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 io_in[21] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
Xinput24 la1_data_in[26] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3460_ _4223_/A _3557_/B vssd1 vssd1 vccd1 vccd1 _3467_/A sky130_fd_sc_hd__or2_2
X_3391_ _4899_/Q _3363_/X _3389_/Y _3390_/X _3325_/X vssd1 vssd1 vccd1 vccd1 _4899_/D
+ sky130_fd_sc_hd__o221a_1
X_5061_ _5099_/CLK _5061_/D vssd1 vssd1 vccd1 vccd1 _5061_/Q sky130_fd_sc_hd__dfxtp_1
X_4012_ _4003_/A _4005_/X _4010_/Y _3943_/A vssd1 vssd1 vccd1 vccd1 _4012_/X sky130_fd_sc_hd__a31o_1
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4914_ _5094_/CLK _4914_/D vssd1 vssd1 vccd1 vccd1 _4914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4845_ _5121_/CLK _4845_/D vssd1 vssd1 vccd1 vccd1 _4845_/Q sky130_fd_sc_hd__dfxtp_1
X_4776_ _4995_/CLK _4776_/D vssd1 vssd1 vccd1 vccd1 _4776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3727_ _5121_/Q _4953_/Q vssd1 vssd1 vccd1 vccd1 _3728_/B sky130_fd_sc_hd__nand2_1
X_3658_ _4022_/A vssd1 vssd1 vccd1 vccd1 _3945_/A sky130_fd_sc_hd__clkbuf_2
X_2609_ _2609_/A _2609_/B vssd1 vssd1 vccd1 vccd1 _2610_/A sky130_fd_sc_hd__and2_1
X_3589_ _3575_/A _3575_/B _3580_/Y _3588_/X vssd1 vssd1 vccd1 vccd1 _3590_/B sky130_fd_sc_hd__a31o_1
X_5259_ _5259_/A _2449_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2960_ _3168_/B _2965_/B vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__nand2_1
X_2891_ _2878_/X _4826_/Q _2888_/X _2890_/X _2876_/X vssd1 vssd1 vccd1 vccd1 _4826_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4630_ _4644_/A _4630_/B vssd1 vssd1 vccd1 vccd1 _4631_/A sky130_fd_sc_hd__and2_1
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4561_ _4892_/Q _5072_/Q _4561_/S vssd1 vssd1 vccd1 vccd1 _4562_/B sky130_fd_sc_hd__mux2_1
X_4492_ _4505_/A _4492_/B vssd1 vssd1 vccd1 vccd1 _4493_/A sky130_fd_sc_hd__and2_1
X_3512_ _4927_/Q _5095_/Q vssd1 vssd1 vccd1 vccd1 _3521_/B sky130_fd_sc_hd__and2_1
X_3443_ _4918_/Q _5086_/Q vssd1 vssd1 vccd1 vccd1 _3445_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3374_ _3371_/X _3372_/Y _3373_/X vssd1 vssd1 vccd1 vccd1 _3374_/X sky130_fd_sc_hd__a21o_1
X_5113_ _5114_/CLK _5113_/D vssd1 vssd1 vccd1 vccd1 _5113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5044_ _5046_/CLK _5044_/D vssd1 vssd1 vccd1 vccd1 _5044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4828_ _4836_/CLK _4828_/D vssd1 vssd1 vccd1 vccd1 _4828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4759_ _4978_/CLK _4759_/D vssd1 vssd1 vccd1 vccd1 _4759_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4989_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3090_ _4874_/Q _5042_/Q vssd1 vssd1 vccd1 vccd1 _3092_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3992_ _3992_/A _4767_/Q vssd1 vssd1 vccd1 vccd1 _3992_/X sky130_fd_sc_hd__or2_1
X_2943_ _2943_/A vssd1 vssd1 vccd1 vccd1 _4839_/D sky130_fd_sc_hd__clkbuf_1
X_2874_ _2862_/X input6/X _2863_/X vssd1 vssd1 vccd1 vccd1 _2874_/X sky130_fd_sc_hd__o21a_1
X_4613_ _4626_/A _4613_/B vssd1 vssd1 vccd1 vccd1 _4614_/A sky130_fd_sc_hd__and2_1
X_4544_ _4544_/A vssd1 vssd1 vccd1 vccd1 _5067_/D sky130_fd_sc_hd__clkbuf_1
X_5166__73 vssd1 vssd1 vccd1 vccd1 _5166__73/HI _5261_/A sky130_fd_sc_hd__conb_1
X_4475_ _4488_/A _4475_/B vssd1 vssd1 vccd1 vccd1 _4476_/A sky130_fd_sc_hd__and2_1
X_3426_ _3424_/Y _3422_/C _3425_/X _3421_/C vssd1 vssd1 vccd1 vccd1 _3426_/X sky130_fd_sc_hd__a22o_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _4907_/Q _5075_/Q vssd1 vssd1 vccd1 vccd1 _3357_/X sky130_fd_sc_hd__xor2_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ _3288_/A vssd1 vssd1 vccd1 vccd1 _3288_/X sky130_fd_sc_hd__clkbuf_2
X_5027_ _5027_/CLK _5027_/D vssd1 vssd1 vccd1 vccd1 _5027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5204__111 vssd1 vssd1 vccd1 vccd1 _5204__111/HI _5312_/A sky130_fd_sc_hd__conb_1
XFILLER_29_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2590_ _2625_/A vssd1 vssd1 vccd1 vccd1 _2604_/S sky130_fd_sc_hd__clkbuf_4
X_4260_ _4284_/A _4256_/B _4252_/A vssd1 vssd1 vccd1 vccd1 _4264_/A sky130_fd_sc_hd__a21oi_1
X_4191_ _5010_/Q _4790_/Q _4191_/C vssd1 vssd1 vccd1 vccd1 _4191_/X sky130_fd_sc_hd__and3_1
X_3211_ _3233_/A _3207_/B _3203_/A vssd1 vssd1 vccd1 vccd1 _3215_/A sky130_fd_sc_hd__a21oi_1
X_3142_ _4880_/Q _5048_/Q vssd1 vssd1 vccd1 vccd1 _3144_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3073_ _3161_/B vssd1 vssd1 vccd1 vccd1 _3074_/A sky130_fd_sc_hd__buf_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3975_ _4985_/Q _4765_/Q vssd1 vssd1 vccd1 vccd1 _3977_/A sky130_fd_sc_hd__nor2_1
X_2926_ _5276_/A _4851_/Q _2968_/B vssd1 vssd1 vccd1 vccd1 _2927_/B sky130_fd_sc_hd__mux2_1
X_2857_ input2/X vssd1 vssd1 vccd1 vccd1 _2889_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2788_ _2919_/A vssd1 vssd1 vccd1 vccd1 _2803_/A sky130_fd_sc_hd__clkbuf_2
X_4527_ _4527_/A vssd1 vssd1 vccd1 vccd1 _5062_/D sky130_fd_sc_hd__clkbuf_1
X_4458_ _4632_/A vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3409_ _4914_/Q _5082_/Q vssd1 vssd1 vccd1 vccd1 _3421_/A sky130_fd_sc_hd__xor2_1
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4389_ _4829_/Q _4817_/Q vssd1 vssd1 vccd1 vccd1 _4389_/Y sky130_fd_sc_hd__nor2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _3754_/A _3754_/B _3759_/Y vssd1 vssd1 vccd1 vccd1 _3765_/A sky130_fd_sc_hd__o21ai_1
X_2711_ _2715_/A _2711_/B vssd1 vssd1 vccd1 vccd1 _2712_/A sky130_fd_sc_hd__and2_1
XFILLER_71_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3691_ _3656_/X _3689_/X _3690_/X _3659_/X vssd1 vssd1 vccd1 vccd1 _4936_/D sky130_fd_sc_hd__o211a_1
X_2642_ _4719_/A vssd1 vssd1 vccd1 vccd1 _2713_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5136__43 vssd1 vssd1 vccd1 vccd1 _5136__43/HI _5231_/A sky130_fd_sc_hd__conb_1
X_2573_ _2625_/A vssd1 vssd1 vccd1 vccd1 _2587_/S sky130_fd_sc_hd__clkbuf_2
X_5292_ _5292_/A _2488_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
X_4312_ _5015_/Q _4259_/X _4310_/X _4311_/Y _4281_/X vssd1 vssd1 vccd1 vccd1 _5015_/D
+ sky130_fd_sc_hd__o221a_1
X_4243_ _4234_/Y _4224_/X _4242_/Y _3360_/X vssd1 vssd1 vccd1 vccd1 _5006_/D sky130_fd_sc_hd__a211oi_1
X_4174_ _4189_/A vssd1 vssd1 vccd1 vccd1 _4174_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3125_ _3138_/A _3109_/B _3115_/A _3137_/A _3124_/Y vssd1 vssd1 vccd1 vccd1 _3125_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_55_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3056_ _4857_/Q _2976_/A _3054_/Y _3055_/X _3037_/X vssd1 vssd1 vccd1 vccd1 _4857_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3958_ _4983_/Q _4763_/Q vssd1 vssd1 vccd1 vccd1 _3959_/B sky130_fd_sc_hd__and2_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3889_ _3883_/A _3882_/B _3887_/Y _3888_/Y vssd1 vssd1 vccd1 vccd1 _3889_/X sky130_fd_sc_hd__a211o_1
X_2909_ _4847_/Q vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4930_ _5121_/CLK _4930_/D vssd1 vssd1 vccd1 vccd1 _4930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4861_ _5040_/CLK _4861_/D vssd1 vssd1 vccd1 vccd1 _4861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3812_ _4964_/Q _4744_/Q vssd1 vssd1 vccd1 vccd1 _3814_/A sky130_fd_sc_hd__nand2_1
X_4792_ _4999_/CLK _4792_/D vssd1 vssd1 vccd1 vccd1 _4792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3743_ _4943_/Q _3664_/A _3741_/X _3742_/Y _3646_/X vssd1 vssd1 vccd1 vccd1 _4943_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3674_ _3672_/X _3673_/Y _3656_/X vssd1 vssd1 vccd1 vccd1 _3674_/Y sky130_fd_sc_hd__a21oi_1
X_2625_ _2625_/A vssd1 vssd1 vccd1 vccd1 _2639_/S sky130_fd_sc_hd__buf_2
X_2556_ _4943_/Q _4735_/Q _2570_/S vssd1 vssd1 vccd1 vccd1 _2557_/B sky130_fd_sc_hd__mux2_1
X_2487_ _2490_/A vssd1 vssd1 vccd1 vccd1 _2487_/Y sky130_fd_sc_hd__inv_2
X_5275_ _5275_/A _2469_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
X_4226_ _5004_/Q _4220_/X _4225_/X _4163_/X vssd1 vssd1 vccd1 vccd1 _5004_/D sky130_fd_sc_hd__o211a_1
X_4157_ _4157_/A _4157_/B vssd1 vssd1 vccd1 vccd1 _4190_/A sky130_fd_sc_hd__nor2_1
XFILLER_28_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3108_ _3094_/A _3094_/B _3099_/Y _3107_/X vssd1 vssd1 vccd1 vccd1 _3109_/B sky130_fd_sc_hd__a31o_2
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4088_ _4999_/Q _4779_/Q vssd1 vssd1 vccd1 vccd1 _4096_/C sky130_fd_sc_hd__or2_1
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_37_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5070_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3039_ _3039_/A _3039_/B _3041_/C vssd1 vssd1 vccd1 vccd1 _3040_/C sky130_fd_sc_hd__and3_1
XFILLER_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput25 la1_data_in[27] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_2
Xinput14 io_in[22] vssd1 vssd1 vccd1 vccd1 _2906_/B sky130_fd_sc_hd__buf_2
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3390_ _3381_/A _3383_/Y _3388_/Y _3373_/X vssd1 vssd1 vccd1 vccd1 _3390_/X sky130_fd_sc_hd__a31o_1
XFILLER_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5060_ _5062_/CLK _5060_/D vssd1 vssd1 vccd1 vccd1 _5060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4011_ _4003_/A _4005_/X _4010_/Y vssd1 vssd1 vccd1 vccd1 _4011_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4913_ _5101_/CLK _4913_/D vssd1 vssd1 vccd1 vccd1 _4913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4844_ _5051_/CLK _4844_/D vssd1 vssd1 vccd1 vccd1 _4844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4775_ _4983_/CLK _4775_/D vssd1 vssd1 vccd1 vccd1 _4775_/Q sky130_fd_sc_hd__dfxtp_1
X_3726_ _5121_/Q _4953_/Q vssd1 vssd1 vccd1 vccd1 _3726_/Y sky130_fd_sc_hd__nor2_1
X_3657_ _3663_/A _3654_/X _3656_/X vssd1 vssd1 vccd1 vccd1 _3657_/X sky130_fd_sc_hd__a21o_1
X_2608_ _4958_/Q _4750_/Q _2622_/S vssd1 vssd1 vccd1 vccd1 _2609_/B sky130_fd_sc_hd__mux2_1
X_3588_ _4934_/Q _5102_/Q _3587_/X _3580_/B vssd1 vssd1 vccd1 vccd1 _3588_/X sky130_fd_sc_hd__a31o_1
X_2539_ _2539_/A vssd1 vssd1 vccd1 vccd1 _2539_/Y sky130_fd_sc_hd__inv_2
X_5258_ _5258_/A _2447_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4209_ _4209_/A _4209_/B vssd1 vssd1 vccd1 vccd1 _4211_/A sky130_fd_sc_hd__or2_1
XFILLER_73_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2890_ _2889_/X input24/X _2883_/X vssd1 vssd1 vccd1 vccd1 _2890_/X sky130_fd_sc_hd__a21bo_1
X_4560_ _4628_/A vssd1 vssd1 vccd1 vccd1 _4575_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4491_ _4872_/Q _5052_/Q _4491_/S vssd1 vssd1 vccd1 vccd1 _4492_/B sky130_fd_sc_hd__mux2_1
X_3511_ _4926_/Q _5094_/Q vssd1 vssd1 vccd1 vccd1 _3520_/A sky130_fd_sc_hd__nand2_1
X_3442_ _4905_/Q _3401_/X _3439_/Y _3440_/X _3441_/X vssd1 vssd1 vccd1 vccd1 _4905_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _3373_/A vssd1 vssd1 vccd1 vccd1 _3373_/X sky130_fd_sc_hd__clkbuf_2
X_5112_ _5117_/CLK _5112_/D vssd1 vssd1 vccd1 vccd1 _5112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5043_ _5046_/CLK _5043_/D vssd1 vssd1 vccd1 vccd1 _5043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4827_ _5040_/CLK _4827_/D vssd1 vssd1 vccd1 vccd1 _4827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4758_ _4978_/CLK _4758_/D vssd1 vssd1 vccd1 vccd1 _4758_/Q sky130_fd_sc_hd__dfxtp_1
X_4689_ _4929_/Q _5109_/Q _4699_/S vssd1 vssd1 vccd1 vccd1 _4690_/B sky130_fd_sc_hd__mux2_1
X_3709_ _3711_/B _3711_/C _3707_/Y _3680_/X vssd1 vssd1 vccd1 vccd1 _3709_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _3992_/A _4767_/Q vssd1 vssd1 vccd1 vccd1 _3991_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2942_ _2951_/A _2942_/B vssd1 vssd1 vccd1 vccd1 _2943_/A sky130_fd_sc_hd__and2_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2873_ _2855_/X _4822_/Q _2871_/X _2872_/X _2869_/X vssd1 vssd1 vccd1 vccd1 _4822_/D
+ sky130_fd_sc_hd__o221a_1
X_4612_ _4907_/Q _5087_/Q _4612_/S vssd1 vssd1 vccd1 vccd1 _4613_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4543_ _4557_/A _4543_/B vssd1 vssd1 vccd1 vccd1 _4544_/A sky130_fd_sc_hd__and2_1
X_4474_ _4867_/Q _5047_/Q _4474_/S vssd1 vssd1 vccd1 vccd1 _4475_/B sky130_fd_sc_hd__mux2_1
X_3425_ _4915_/Q _5083_/Q _5082_/Q _4914_/Q vssd1 vssd1 vccd1 vccd1 _3425_/X sky130_fd_sc_hd__a22o_1
X_5181__88 vssd1 vssd1 vccd1 vccd1 _5181__88/HI _5289_/A sky130_fd_sc_hd__conb_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _3336_/A _3338_/Y _3343_/B _3351_/A _3341_/Y vssd1 vssd1 vccd1 vccd1 _3356_/X
+ sky130_fd_sc_hd__a311o_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3287_/A _3287_/B vssd1 vssd1 vccd1 vccd1 _3287_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5026_/CLK _5026_/D vssd1 vssd1 vccd1 vccd1 _5026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4190_ _4190_/A _4190_/B _4190_/C vssd1 vssd1 vccd1 vccd1 _4190_/X sky130_fd_sc_hd__and3_1
X_3210_ _3176_/X _3207_/X _3208_/X _3209_/X vssd1 vssd1 vccd1 vccd1 _4876_/D sky130_fd_sc_hd__o211a_1
XFILLER_79_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3141_ _3109_/B _3138_/X _3140_/X vssd1 vssd1 vccd1 vccd1 _3146_/A sky130_fd_sc_hd__a21o_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3072_ _4219_/A _3175_/A vssd1 vssd1 vccd1 vccd1 _3161_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3974_ _3971_/A _3971_/B _3966_/A vssd1 vssd1 vccd1 vccd1 _3978_/A sky130_fd_sc_hd__a21oi_1
X_2925_ _2925_/A vssd1 vssd1 vccd1 vccd1 _4834_/D sky130_fd_sc_hd__clkbuf_1
X_2856_ _2856_/A vssd1 vssd1 vccd1 vccd1 _2905_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2787_ _4646_/A vssd1 vssd1 vccd1 vccd1 _2919_/A sky130_fd_sc_hd__clkbuf_2
X_4526_ _4539_/A _4526_/B vssd1 vssd1 vccd1 vccd1 _4527_/A sky130_fd_sc_hd__and2_1
X_4457_ _4457_/A vssd1 vssd1 vccd1 vccd1 _5042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3408_ _4901_/Q _3401_/X _3406_/Y _3407_/X _3325_/X vssd1 vssd1 vccd1 vccd1 _4901_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4388_ _5024_/Q _4315_/X _4387_/X _2869_/X vssd1 vssd1 vccd1 vccd1 _5024_/D sky130_fd_sc_hd__o211a_1
X_3339_ _3337_/X _3338_/Y _3288_/X vssd1 vssd1 vccd1 vccd1 _3339_/X sky130_fd_sc_hd__a21o_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ _5010_/CLK _5009_/D vssd1 vssd1 vccd1 vccd1 _5009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2710_ _3992_/A _4779_/Q _2710_/S vssd1 vssd1 vccd1 vccd1 _2711_/B sky130_fd_sc_hd__mux2_1
X_3690_ _4936_/Q _3737_/B vssd1 vssd1 vccd1 vccd1 _3690_/X sky130_fd_sc_hd__or2_1
X_2641_ _2641_/A vssd1 vssd1 vccd1 vccd1 _4759_/D sky130_fd_sc_hd__clkbuf_1
X_2572_ _2572_/A vssd1 vssd1 vccd1 vccd1 _4739_/D sky130_fd_sc_hd__clkbuf_1
X_5291_ _5291_/A _2487_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
X_4311_ _4303_/B _4308_/Y _4309_/Y _4259_/X vssd1 vssd1 vccd1 vccd1 _4311_/Y sky130_fd_sc_hd__o31ai_1
X_4242_ _4240_/X _4241_/Y _4224_/X vssd1 vssd1 vccd1 vccd1 _4242_/Y sky130_fd_sc_hd__a21oi_1
X_5151__58 vssd1 vssd1 vccd1 vccd1 _5151__58/HI _5246_/A sky130_fd_sc_hd__conb_1
X_4173_ _5010_/Q _4790_/Q vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__xor2_1
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3124_ _3123_/Y _3115_/B _3121_/Y vssd1 vssd1 vccd1 vccd1 _3124_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3055_ _3046_/A _3048_/Y _3053_/X _2988_/A vssd1 vssd1 vccd1 vccd1 _3055_/X sky130_fd_sc_hd__a31o_1
XFILLER_48_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3957_ _4983_/Q _4763_/Q vssd1 vssd1 vccd1 vccd1 _3959_/A sky130_fd_sc_hd__nor2_1
X_2908_ _2855_/X _4831_/Q _2557_/A _2907_/X vssd1 vssd1 vccd1 vccd1 _4831_/D sky130_fd_sc_hd__o211a_1
X_3888_ _4973_/Q _4753_/Q vssd1 vssd1 vccd1 vccd1 _3888_/Y sky130_fd_sc_hd__nor2_1
X_2839_ _2839_/A vssd1 vssd1 vccd1 vccd1 _4815_/D sky130_fd_sc_hd__clkbuf_1
X_4509_ _4522_/A _4509_/B vssd1 vssd1 vccd1 vccd1 _4510_/A sky130_fd_sc_hd__and2_1
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5010_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _5050_/CLK _4860_/D vssd1 vssd1 vccd1 vccd1 _4860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3811_ _3781_/B _3806_/X _3810_/X vssd1 vssd1 vccd1 vccd1 _3816_/A sky130_fd_sc_hd__a21o_1
X_4791_ _4999_/CLK _4791_/D vssd1 vssd1 vccd1 vccd1 _4791_/Q sky130_fd_sc_hd__dfxtp_1
X_3742_ _3734_/B _3739_/Y _3740_/Y _3737_/B vssd1 vssd1 vccd1 vccd1 _3742_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3673_ _3673_/A _3673_/B vssd1 vssd1 vccd1 vccd1 _3673_/Y sky130_fd_sc_hd__nand2_1
X_2624_ _2624_/A vssd1 vssd1 vccd1 vccd1 _4754_/D sky130_fd_sc_hd__clkbuf_1
X_2555_ _2625_/A vssd1 vssd1 vccd1 vccd1 _2570_/S sky130_fd_sc_hd__clkbuf_4
X_2486_ _2490_/A vssd1 vssd1 vccd1 vccd1 _2486_/Y sky130_fd_sc_hd__inv_2
X_5274_ _5274_/A _2468_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
X_4225_ _4221_/X _4229_/A _4224_/X vssd1 vssd1 vccd1 vccd1 _4225_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4156_ _5008_/Q _4788_/Q vssd1 vssd1 vccd1 vccd1 _4157_/B sky130_fd_sc_hd__nor2_1
X_3107_ _4874_/Q _5042_/Q _3106_/X _3099_/B vssd1 vssd1 vccd1 vccd1 _3107_/X sky130_fd_sc_hd__a31o_1
X_4087_ _4999_/Q _4779_/Q vssd1 vssd1 vccd1 vccd1 _4092_/B sky130_fd_sc_hd__nand2_1
X_3038_ _4855_/Q _2976_/A _3035_/Y _3036_/X _3037_/X vssd1 vssd1 vccd1 vccd1 _4855_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4989_ _4989_/CLK _4989_/D vssd1 vssd1 vccd1 vccd1 _4989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput26 la1_data_in[28] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput15 io_in[8] vssd1 vssd1 vccd1 vccd1 _3168_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4010_ _4010_/A _4010_/B vssd1 vssd1 vccd1 vccd1 _4010_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ _5091_/CLK _4912_/D vssd1 vssd1 vccd1 vccd1 _4912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4843_ _5050_/CLK _4843_/D vssd1 vssd1 vccd1 vccd1 _5284_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4774_ _4981_/CLK _4774_/D vssd1 vssd1 vccd1 vccd1 _4774_/Q sky130_fd_sc_hd__dfxtp_1
X_3725_ _4940_/Q _3652_/X _3723_/X _3724_/X vssd1 vssd1 vccd1 vccd1 _4940_/D sky130_fd_sc_hd__o211a_1
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3656_ _3680_/A vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__buf_2
X_2607_ _2625_/A vssd1 vssd1 vccd1 vccd1 _2622_/S sky130_fd_sc_hd__buf_2
X_3587_ _4935_/Q _5103_/Q vssd1 vssd1 vccd1 vccd1 _3587_/X sky130_fd_sc_hd__or2_1
X_2538_ _2539_/A vssd1 vssd1 vccd1 vccd1 _2538_/Y sky130_fd_sc_hd__inv_2
X_5257_ _5257_/A _2446_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4208_ _5014_/Q _4794_/Q vssd1 vssd1 vccd1 vccd1 _4209_/B sky130_fd_sc_hd__and2_1
X_2469_ _2472_/A vssd1 vssd1 vccd1 vccd1 _2469_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4139_ _4994_/Q vssd1 vssd1 vccd1 vccd1 _4139_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5187__94 vssd1 vssd1 vccd1 vccd1 _5187__94/HI _5295_/A sky130_fd_sc_hd__conb_1
XFILLER_78_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3510_ _4914_/Q _3457_/X _3509_/X _3503_/X vssd1 vssd1 vccd1 vccd1 _4914_/D sky130_fd_sc_hd__o211a_1
X_4490_ _4541_/A vssd1 vssd1 vccd1 vccd1 _4505_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3441_ _3551_/A vssd1 vssd1 vccd1 vccd1 _3441_/X sky130_fd_sc_hd__clkbuf_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3372_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3372_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5111_ _5121_/CLK _5111_/D vssd1 vssd1 vccd1 vccd1 _5111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5042_ _5046_/CLK _5042_/D vssd1 vssd1 vccd1 vccd1 _5042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4826_ _5040_/CLK _4826_/D vssd1 vssd1 vccd1 vccd1 _4826_/Q sky130_fd_sc_hd__dfxtp_1
X_4757_ _4978_/CLK _4757_/D vssd1 vssd1 vccd1 vccd1 _4757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4688_ _4688_/A vssd1 vssd1 vccd1 vccd1 _5108_/D sky130_fd_sc_hd__clkbuf_1
X_3708_ _3711_/B _3711_/C _3707_/Y vssd1 vssd1 vccd1 vccd1 _3708_/Y sky130_fd_sc_hd__a21oi_1
X_3639_ _4930_/Q _3639_/B vssd1 vssd1 vccd1 vccd1 _3639_/X sky130_fd_sc_hd__or2_1
X_5309_ _5309_/A _2509_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4752_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3990_ _3995_/A _3983_/X _3996_/B _3996_/C vssd1 vssd1 vccd1 vccd1 _3990_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2941_ _5280_/A _4855_/Q _2944_/S vssd1 vssd1 vccd1 vccd1 _2942_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ _4628_/A vssd1 vssd1 vccd1 vccd1 _4626_/A sky130_fd_sc_hd__clkbuf_2
X_2872_ _2865_/X input20/X _2878_/A vssd1 vssd1 vccd1 vccd1 _2872_/X sky130_fd_sc_hd__a21bo_1
X_4542_ _4887_/Q _5067_/Q _4542_/S vssd1 vssd1 vccd1 vccd1 _4543_/B sky130_fd_sc_hd__mux2_1
X_4473_ _4541_/A vssd1 vssd1 vccd1 vccd1 _4488_/A sky130_fd_sc_hd__clkbuf_2
X_3424_ _3423_/Y _3405_/B _3403_/Y vssd1 vssd1 vccd1 vccd1 _3424_/Y sky130_fd_sc_hd__a21oi_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _4895_/Q vssd1 vssd1 vccd1 vccd1 _3355_/Y sky130_fd_sc_hd__inv_2
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3287_/A _3287_/B vssd1 vssd1 vccd1 vccd1 _3286_/X sky130_fd_sc_hd__or2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5027_/CLK _5025_/D vssd1 vssd1 vccd1 vccd1 _5025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4809_ _5018_/CLK _4809_/D vssd1 vssd1 vccd1 vccd1 _4809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5157__64 vssd1 vssd1 vccd1 vccd1 _5157__64/HI _5252_/A sky130_fd_sc_hd__conb_1
XFILLER_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3140_ _4879_/Q _5047_/Q _3124_/Y _3138_/C _3139_/X vssd1 vssd1 vccd1 vccd1 _3140_/X
+ sky130_fd_sc_hd__a221o_1
X_3071_ _4223_/A vssd1 vssd1 vccd1 vccd1 _4219_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ _4972_/Q _3933_/X _3972_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _4972_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2924_ _2934_/A _2924_/B vssd1 vssd1 vccd1 vccd1 _2925_/A sky130_fd_sc_hd__and2_1
X_2855_ _2855_/A vssd1 vssd1 vccd1 vccd1 _2855_/X sky130_fd_sc_hd__clkbuf_2
X_4525_ _4882_/Q _5062_/Q _4525_/S vssd1 vssd1 vccd1 vccd1 _4526_/B sky130_fd_sc_hd__mux2_1
X_2786_ _3133_/A vssd1 vssd1 vccd1 vccd1 _4646_/A sky130_fd_sc_hd__buf_4
X_4456_ _4470_/A _4456_/B vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__and2_1
X_3407_ _3406_/A _3422_/B _3373_/X vssd1 vssd1 vccd1 vccd1 _3407_/X sky130_fd_sc_hd__a21o_1
X_4387_ _4385_/X _4386_/Y _4326_/X vssd1 vssd1 vccd1 vccd1 _4387_/X sky130_fd_sc_hd__a21o_1
X_3338_ _3338_/A _3338_/B vssd1 vssd1 vccd1 vccd1 _3338_/Y sky130_fd_sc_hd__nand2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3269_ _4896_/Q _5064_/Q vssd1 vssd1 vccd1 vccd1 _3269_/X sky130_fd_sc_hd__or2_1
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _5010_/CLK _5008_/D vssd1 vssd1 vccd1 vccd1 _5008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2640_ _2645_/A _2640_/B vssd1 vssd1 vccd1 vccd1 _2641_/A sky130_fd_sc_hd__and2_1
X_2571_ _2575_/A _2571_/B vssd1 vssd1 vccd1 vccd1 _2572_/A sky130_fd_sc_hd__and2_1
X_5290_ _5290_/A _2486_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
X_4310_ _4303_/B _4308_/Y _4309_/Y vssd1 vssd1 vccd1 vccd1 _4310_/X sky130_fd_sc_hd__o21a_1
X_4241_ _4241_/A _4241_/B vssd1 vssd1 vccd1 vccd1 _4241_/Y sky130_fd_sc_hd__nand2_1
X_4172_ _4997_/Q _4165_/X _4170_/Y _4171_/X _4076_/X vssd1 vssd1 vccd1 vccd1 _4997_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3123_ _4876_/Q _5044_/Q vssd1 vssd1 vccd1 vccd1 _3123_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3054_ _3046_/A _3048_/Y _3053_/X vssd1 vssd1 vccd1 vccd1 _3054_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3956_ _3947_/Y _3937_/X _3955_/Y _3360_/X vssd1 vssd1 vccd1 vccd1 _4970_/D sky130_fd_sc_hd__a211oi_1
X_2907_ _2905_/X _2906_/X _2855_/A vssd1 vssd1 vccd1 vccd1 _2907_/X sky130_fd_sc_hd__a21bo_1
X_3887_ _3901_/A vssd1 vssd1 vccd1 vccd1 _3887_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2838_ _2838_/A _2838_/B vssd1 vssd1 vccd1 vccd1 _2839_/A sky130_fd_sc_hd__and2_1
X_2769_ _2769_/A vssd1 vssd1 vccd1 vccd1 _2784_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4508_ _4877_/Q _5057_/Q _4508_/S vssd1 vssd1 vccd1 vccd1 _4509_/B sky130_fd_sc_hd__mux2_1
X_5127__34 vssd1 vssd1 vccd1 vccd1 _5127__34/HI _5222_/A sky130_fd_sc_hd__conb_1
X_4439_ _4452_/A _4439_/B vssd1 vssd1 vccd1 vccd1 _4440_/A sky130_fd_sc_hd__and2_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4790_ _4999_/CLK _4790_/D vssd1 vssd1 vccd1 vccd1 _4790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3810_ _3808_/Y _3806_/C _3809_/X _3805_/C vssd1 vssd1 vccd1 vccd1 _3810_/X sky130_fd_sc_hd__a22o_1
X_3741_ _3734_/B _3739_/Y _3740_/Y vssd1 vssd1 vccd1 vccd1 _3741_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3672_ _3673_/A _3673_/B vssd1 vssd1 vccd1 vccd1 _3672_/X sky130_fd_sc_hd__or2_1
X_2623_ _2627_/A _2623_/B vssd1 vssd1 vccd1 vccd1 _2624_/A sky130_fd_sc_hd__and2_1
X_2554_ _4719_/A vssd1 vssd1 vccd1 vccd1 _2625_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2485_ _2485_/A vssd1 vssd1 vccd1 vccd1 _2490_/A sky130_fd_sc_hd__buf_12
X_5273_ _5273_/A _2466_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
X_4224_ _4230_/A vssd1 vssd1 vccd1 vccd1 _4224_/X sky130_fd_sc_hd__clkbuf_2
X_4155_ _5008_/Q _4788_/Q vssd1 vssd1 vccd1 vccd1 _4157_/A sky130_fd_sc_hd__and2_1
X_3106_ _4875_/Q _5043_/Q vssd1 vssd1 vccd1 vccd1 _3106_/X sky130_fd_sc_hd__or2_1
X_4086_ _4086_/A _4086_/B vssd1 vssd1 vccd1 vccd1 _4086_/X sky130_fd_sc_hd__or2_1
X_3037_ _3037_/A vssd1 vssd1 vccd1 vccd1 _3037_/X sky130_fd_sc_hd__buf_2
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4988_ _4989_/CLK _4988_/D vssd1 vssd1 vccd1 vccd1 _4988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3939_ _4968_/Q _3933_/X _3938_/X _3876_/X vssd1 vssd1 vccd1 vccd1 _4968_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_46_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5046_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 io_in[9] vssd1 vssd1 vccd1 vccd1 _2856_/A sky130_fd_sc_hd__clkbuf_2
Xinput27 la1_data_in[29] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ _5101_/CLK _4911_/D vssd1 vssd1 vccd1 vccd1 _4911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4842_ _5041_/CLK _4842_/D vssd1 vssd1 vccd1 vccd1 _5283_/A sky130_fd_sc_hd__dfxtp_1
X_4773_ _4983_/CLK _4773_/D vssd1 vssd1 vccd1 vccd1 _4773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3724_ _3945_/A vssd1 vssd1 vccd1 vccd1 _3724_/X sky130_fd_sc_hd__buf_2
X_3655_ _4032_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _3680_/A sky130_fd_sc_hd__or2_1
X_2606_ _2606_/A vssd1 vssd1 vccd1 vccd1 _4749_/D sky130_fd_sc_hd__clkbuf_1
X_3586_ _3586_/A _3586_/B vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__nor2_1
X_2537_ _2539_/A vssd1 vssd1 vccd1 vccd1 _2537_/Y sky130_fd_sc_hd__inv_2
X_5325_ _5325_/A _2529_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
X_5256_ _5256_/A _2445_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
X_2468_ _2472_/A vssd1 vssd1 vccd1 vccd1 _2468_/Y sky130_fd_sc_hd__inv_2
X_4207_ _5014_/Q _4794_/Q vssd1 vssd1 vccd1 vccd1 _4209_/A sky130_fd_sc_hd__nor2_1
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4138_ _4993_/Q _4126_/X _4137_/X _4082_/X vssd1 vssd1 vccd1 vccd1 _4993_/D sky130_fd_sc_hd__o211a_1
X_4069_ _4038_/X _4067_/X _4068_/X _4023_/X vssd1 vssd1 vccd1 vccd1 _4984_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3440_ _3430_/A _3432_/Y _3438_/X _3373_/A vssd1 vssd1 vccd1 vccd1 _3440_/X sky130_fd_sc_hd__a31o_1
X_3371_ _3372_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3371_/X sky130_fd_sc_hd__or2_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5110_ _5121_/CLK _5110_/D vssd1 vssd1 vccd1 vccd1 _5110_/Q sky130_fd_sc_hd__dfxtp_1
X_5041_ _5041_/CLK _5041_/D vssd1 vssd1 vccd1 vccd1 _5041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_80_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4825_ _5050_/CLK _4825_/D vssd1 vssd1 vccd1 vccd1 _4825_/Q sky130_fd_sc_hd__dfxtp_1
X_4756_ _4972_/CLK _4756_/D vssd1 vssd1 vccd1 vccd1 _4756_/Q sky130_fd_sc_hd__dfxtp_1
X_4687_ _4696_/A _4687_/B vssd1 vssd1 vccd1 vccd1 _4688_/A sky130_fd_sc_hd__and2_1
X_3707_ _5118_/Q _4950_/Q _3711_/A _3702_/B vssd1 vssd1 vccd1 vccd1 _3707_/Y sky130_fd_sc_hd__a22oi_1
X_3638_ _3638_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _3638_/X sky130_fd_sc_hd__xor2_1
X_3569_ _4933_/Q _5101_/Q vssd1 vssd1 vccd1 vccd1 _3569_/Y sky130_fd_sc_hd__nand2_1
X_5308_ _5308_/A _2508_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
X_5239_ _5239_/A _2537_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2940_ _2940_/A vssd1 vssd1 vccd1 vccd1 _4838_/D sky130_fd_sc_hd__clkbuf_1
X_2871_ _2862_/X input5/X _2863_/X vssd1 vssd1 vccd1 vccd1 _2871_/X sky130_fd_sc_hd__o21a_1
X_4610_ _4610_/A vssd1 vssd1 vccd1 vccd1 _5086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4541_ _4541_/A vssd1 vssd1 vccd1 vccd1 _4557_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4472_ _4646_/A vssd1 vssd1 vccd1 vccd1 _4541_/A sky130_fd_sc_hd__clkbuf_2
X_3423_ _4912_/Q _5080_/Q vssd1 vssd1 vccd1 vccd1 _3423_/Y sky130_fd_sc_hd__nand2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3272_/X _3351_/X _3352_/X _3353_/X vssd1 vssd1 vccd1 vccd1 _4894_/D sky130_fd_sc_hd__o211a_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3285_/A _3285_/B vssd1 vssd1 vccd1 vccd1 _3287_/B sky130_fd_sc_hd__and2_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5026_/CLK _5024_/D vssd1 vssd1 vccd1 vccd1 _5024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4808_ _5018_/CLK _4808_/D vssd1 vssd1 vccd1 vccd1 _4808_/Q sky130_fd_sc_hd__dfxtp_1
X_4739_ _4948_/CLK _4739_/D vssd1 vssd1 vccd1 vccd1 _4739_/Q sky130_fd_sc_hd__dfxtp_1
X_5172__79 vssd1 vssd1 vccd1 vccd1 _5172__79/HI _5267_/A sky130_fd_sc_hd__conb_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5211__118 vssd1 vssd1 vccd1 vccd1 _5211__118/HI _5319_/A sky130_fd_sc_hd__conb_1
XFILLER_5_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3070_ _3168_/A _4845_/Q _4844_/Q vssd1 vssd1 vccd1 vccd1 _4223_/A sky130_fd_sc_hd__or3b_4
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3972_ _3970_/Y _3971_/X _3943_/X vssd1 vssd1 vccd1 vccd1 _3972_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2923_ _5275_/A _4850_/Q _2968_/B vssd1 vssd1 vccd1 vccd1 _2924_/B sky130_fd_sc_hd__mux2_1
X_2854_ _2958_/B vssd1 vssd1 vccd1 vccd1 _2855_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2785_ _2785_/A vssd1 vssd1 vccd1 vccd1 _4800_/D sky130_fd_sc_hd__clkbuf_1
X_4524_ _4541_/A vssd1 vssd1 vccd1 vccd1 _4539_/A sky130_fd_sc_hd__clkbuf_2
X_4455_ _4862_/Q _5042_/Q _4455_/S vssd1 vssd1 vccd1 vccd1 _4456_/B sky130_fd_sc_hd__mux2_1
X_3406_ _3406_/A _3422_/B vssd1 vssd1 vccd1 vccd1 _3406_/Y sky130_fd_sc_hd__nor2_1
X_4386_ _4386_/A _4386_/B vssd1 vssd1 vccd1 vccd1 _4386_/Y sky130_fd_sc_hd__nand2_2
X_3337_ _3338_/A _3338_/B vssd1 vssd1 vccd1 vccd1 _3337_/X sky130_fd_sc_hd__or2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _3277_/A vssd1 vssd1 vccd1 vccd1 _3268_/X sky130_fd_sc_hd__clkbuf_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3199_ _3189_/A _3192_/B _3197_/Y _3182_/X vssd1 vssd1 vccd1 vccd1 _3199_/X sky130_fd_sc_hd__a31o_1
X_5007_ _5026_/CLK _5007_/D vssd1 vssd1 vccd1 vccd1 _5007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2570_ _4947_/Q _4739_/Q _2570_/S vssd1 vssd1 vccd1 vccd1 _2571_/B sky130_fd_sc_hd__mux2_1
XFILLER_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4240_ _4241_/A _4241_/B vssd1 vssd1 vccd1 vccd1 _4240_/X sky130_fd_sc_hd__or2_1
X_4171_ _4170_/A _4190_/B _4136_/X vssd1 vssd1 vccd1 vccd1 _4171_/X sky130_fd_sc_hd__a21o_1
X_3122_ _3116_/A _3115_/B _3120_/Y _3121_/Y vssd1 vssd1 vccd1 vccd1 _3122_/X sky130_fd_sc_hd__a211o_1
X_3053_ _3051_/Y _3053_/B vssd1 vssd1 vccd1 vccd1 _3053_/X sky130_fd_sc_hd__and2b_1
XFILLER_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3955_ _3953_/X _3954_/Y _3937_/X vssd1 vssd1 vccd1 vccd1 _3955_/Y sky130_fd_sc_hd__a21oi_1
X_2906_ input2/X _2906_/B _2856_/A vssd1 vssd1 vccd1 vccd1 _2906_/X sky130_fd_sc_hd__or3b_1
X_3886_ _4974_/Q _4754_/Q vssd1 vssd1 vccd1 vccd1 _3901_/A sky130_fd_sc_hd__xor2_1
X_2837_ _5023_/Q _4815_/Q _2850_/S vssd1 vssd1 vccd1 vccd1 _2838_/B sky130_fd_sc_hd__mux2_1
X_2768_ _2768_/A vssd1 vssd1 vccd1 vccd1 _4795_/D sky130_fd_sc_hd__clkbuf_1
X_2699_ _2769_/A vssd1 vssd1 vccd1 vccd1 _2715_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4507_ _4541_/A vssd1 vssd1 vccd1 vccd1 _4522_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4438_ _4857_/Q _5037_/Q _4438_/S vssd1 vssd1 vccd1 vccd1 _4439_/B sky130_fd_sc_hd__mux2_1
X_5142__49 vssd1 vssd1 vccd1 vccd1 _5142__49/HI _5237_/A sky130_fd_sc_hd__conb_1
X_4369_ _4369_/A _4369_/B vssd1 vssd1 vccd1 vccd1 _4369_/X sky130_fd_sc_hd__or2_1
XFILLER_58_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5217__124 vssd1 vssd1 vccd1 vccd1 _5217__124/HI _5325_/A sky130_fd_sc_hd__conb_1
X_3740_ _4955_/Q _4735_/Q vssd1 vssd1 vccd1 vccd1 _3740_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3671_ _3671_/A _3671_/B vssd1 vssd1 vccd1 vccd1 _3673_/B sky130_fd_sc_hd__and2_1
X_2622_ _4962_/Q _4754_/Q _2622_/S vssd1 vssd1 vccd1 vccd1 _2623_/B sky130_fd_sc_hd__mux2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2553_ _4632_/A vssd1 vssd1 vccd1 vccd1 _4719_/A sky130_fd_sc_hd__buf_2
X_5272_ _5272_/A _2465_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
X_2484_ _2484_/A vssd1 vssd1 vccd1 vccd1 _2484_/Y sky130_fd_sc_hd__inv_2
X_4223_ _4223_/A _4223_/B vssd1 vssd1 vccd1 vccd1 _4230_/A sky130_fd_sc_hd__or2_2
X_4154_ _4995_/Q _4126_/X _4152_/Y _4153_/X _4076_/X vssd1 vssd1 vccd1 vccd1 _4995_/D
+ sky130_fd_sc_hd__o221a_1
X_4085_ _4092_/A vssd1 vssd1 vccd1 vccd1 _4086_/A sky130_fd_sc_hd__clkinv_2
X_3105_ _3105_/A _3105_/B vssd1 vssd1 vccd1 vccd1 _3138_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3036_ _3032_/Y _3026_/X _3039_/B _3041_/C _2988_/A vssd1 vssd1 vccd1 vccd1 _3036_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4987_ _4989_/CLK _4987_/D vssd1 vssd1 vccd1 vccd1 _4987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3938_ _3934_/X _3942_/A _3937_/X vssd1 vssd1 vccd1 vccd1 _3938_/X sky130_fd_sc_hd__a21o_1
X_3869_ _4972_/Q _4752_/Q vssd1 vssd1 vccd1 vccd1 _3870_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5122_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 la1_data_in[0] vssd1 vssd1 vccd1 vccd1 _5285_/A sky130_fd_sc_hd__buf_6
Xinput28 la1_data_in[30] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4910_ _5101_/CLK _4910_/D vssd1 vssd1 vccd1 vccd1 _4910_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4841_ _5040_/CLK _4841_/D vssd1 vssd1 vccd1 vccd1 _5282_/A sky130_fd_sc_hd__dfxtp_1
X_4772_ _4989_/CLK _4772_/D vssd1 vssd1 vccd1 vccd1 _4772_/Q sky130_fd_sc_hd__dfxtp_1
X_3723_ _3721_/X _3722_/Y _3680_/X vssd1 vssd1 vccd1 vccd1 _3723_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3654_ _5112_/Q _4944_/Q vssd1 vssd1 vccd1 vccd1 _3654_/X sky130_fd_sc_hd__or2_1
X_2605_ _2609_/A _2605_/B vssd1 vssd1 vccd1 vccd1 _2606_/A sky130_fd_sc_hd__and2_1
X_3585_ _4936_/Q _5104_/Q vssd1 vssd1 vccd1 vccd1 _3586_/B sky130_fd_sc_hd__nor2_1
X_2536_ _2539_/A vssd1 vssd1 vccd1 vccd1 _2536_/Y sky130_fd_sc_hd__inv_2
X_5324_ _5324_/A _2527_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
X_5255_ _5255_/A _2444_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
X_2467_ _2485_/A vssd1 vssd1 vccd1 vccd1 _2472_/A sky130_fd_sc_hd__clkbuf_4
X_4206_ _5001_/Q _4165_/X _4204_/Y _4205_/X _4187_/X vssd1 vssd1 vccd1 vccd1 _5001_/D
+ sky130_fd_sc_hd__o221a_1
X_4137_ _4134_/X _4135_/Y _4136_/X vssd1 vssd1 vccd1 vccd1 _4137_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4068_ _4984_/Q _4117_/B vssd1 vssd1 vccd1 vccd1 _4068_/X sky130_fd_sc_hd__or2_1
X_3019_ _3019_/A _3019_/B vssd1 vssd1 vccd1 vccd1 _3040_/B sky130_fd_sc_hd__and2_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5178__85 vssd1 vssd1 vccd1 vccd1 _5178__85/HI _5286_/A sky130_fd_sc_hd__conb_1
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3370_ _4909_/Q _5077_/Q vssd1 vssd1 vccd1 vccd1 _3372_/B sky130_fd_sc_hd__xnor2_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/CLK _5040_/D vssd1 vssd1 vccd1 vccd1 _5040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4824_ _5050_/CLK _4824_/D vssd1 vssd1 vccd1 vccd1 _4824_/Q sky130_fd_sc_hd__dfxtp_1
X_4755_ _4972_/CLK _4755_/D vssd1 vssd1 vccd1 vccd1 _4755_/Q sky130_fd_sc_hd__dfxtp_1
X_3706_ _5119_/Q _4951_/Q vssd1 vssd1 vccd1 vccd1 _3711_/C sky130_fd_sc_hd__or2_1
X_4686_ _4928_/Q _5108_/Q _4699_/S vssd1 vssd1 vccd1 vccd1 _4687_/B sky130_fd_sc_hd__mux2_1
X_3637_ _3623_/A _3625_/Y _3630_/B _3628_/Y vssd1 vssd1 vccd1 vccd1 _3638_/B sky130_fd_sc_hd__a31o_1
X_3568_ _4922_/Q vssd1 vssd1 vccd1 vccd1 _3568_/Y sky130_fd_sc_hd__inv_2
X_5307_ _5307_/A _2507_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
X_2519_ _2521_/A vssd1 vssd1 vccd1 vccd1 _2519_/Y sky130_fd_sc_hd__inv_2
X_3499_ _4925_/Q _5093_/Q vssd1 vssd1 vccd1 vccd1 _3499_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5238_ _5238_/A _2535_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5103_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2870_ _2855_/X _4821_/Q _2864_/X _2867_/X _2869_/X vssd1 vssd1 vccd1 vccd1 _4821_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _4540_/A vssd1 vssd1 vccd1 vccd1 _5066_/D sky130_fd_sc_hd__clkbuf_1
X_4471_ _4471_/A vssd1 vssd1 vccd1 vccd1 _5046_/D sky130_fd_sc_hd__clkbuf_1
X_3422_ _3422_/A _3422_/B _3422_/C vssd1 vssd1 vccd1 vccd1 _3422_/X sky130_fd_sc_hd__and3_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3566_/A vssd1 vssd1 vccd1 vccd1 _3353_/X sky130_fd_sc_hd__buf_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _4898_/Q _5066_/Q vssd1 vssd1 vccd1 vccd1 _3285_/B sky130_fd_sc_hd__or2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5026_/CLK _5023_/D vssd1 vssd1 vccd1 vccd1 _5023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4807_ _5015_/CLK _4807_/D vssd1 vssd1 vccd1 vccd1 _4807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2999_ _2997_/X _2998_/Y _2980_/X vssd1 vssd1 vccd1 vccd1 _2999_/Y sky130_fd_sc_hd__a21oi_1
X_4738_ _4948_/CLK _4738_/D vssd1 vssd1 vccd1 vccd1 _4738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4669_ _4923_/Q _5103_/Q _4682_/S vssd1 vssd1 vccd1 vccd1 _4670_/B sky130_fd_sc_hd__mux2_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5148__55 vssd1 vssd1 vccd1 vccd1 _5148__55/HI _5243_/A sky130_fd_sc_hd__conb_1
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3971_ _3971_/A _3971_/B vssd1 vssd1 vccd1 vccd1 _3971_/X sky130_fd_sc_hd__or2_1
X_2922_ _2922_/A vssd1 vssd1 vccd1 vccd1 _4833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2853_ _4719_/A vssd1 vssd1 vccd1 vccd1 _2958_/B sky130_fd_sc_hd__clkbuf_2
X_2784_ _2784_/A _2784_/B vssd1 vssd1 vccd1 vccd1 _2785_/A sky130_fd_sc_hd__and2_1
X_4523_ _4523_/A vssd1 vssd1 vccd1 vccd1 _5061_/D sky130_fd_sc_hd__clkbuf_1
X_4454_ _4454_/A vssd1 vssd1 vccd1 vccd1 _4470_/A sky130_fd_sc_hd__clkbuf_2
X_3405_ _3403_/Y _3405_/B vssd1 vssd1 vccd1 vccd1 _3422_/B sky130_fd_sc_hd__and2b_1
X_4385_ _4386_/A _4386_/B vssd1 vssd1 vccd1 vccd1 _4385_/X sky130_fd_sc_hd__or2_1
X_3336_ _3336_/A _3336_/B vssd1 vssd1 vccd1 vccd1 _3338_/B sky130_fd_sc_hd__and2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3267_ _3352_/B vssd1 vssd1 vccd1 vccd1 _3277_/A sky130_fd_sc_hd__clkbuf_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5026_/CLK _5006_/D vssd1 vssd1 vccd1 vccd1 _5006_/Q sky130_fd_sc_hd__dfxtp_1
X_3198_ _3189_/A _3192_/B _3197_/Y vssd1 vssd1 vccd1 vccd1 _3198_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _4170_/A _4190_/B vssd1 vssd1 vccd1 vccd1 _4170_/Y sky130_fd_sc_hd__nor2_1
X_3121_ _4877_/Q _5045_/Q vssd1 vssd1 vccd1 vccd1 _3121_/Y sky130_fd_sc_hd__nor2_1
X_3052_ _4869_/Q _5037_/Q vssd1 vssd1 vccd1 vccd1 _3053_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3954_ _3954_/A _3954_/B vssd1 vssd1 vccd1 vccd1 _3954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3885_ _4961_/Q _3878_/X _3883_/Y _3884_/X _3866_/X vssd1 vssd1 vccd1 vccd1 _4961_/D
+ sky130_fd_sc_hd__o221a_1
X_2905_ _2905_/A _2905_/B input2/X vssd1 vssd1 vccd1 vccd1 _2905_/X sky130_fd_sc_hd__or3b_1
X_2836_ _4441_/A vssd1 vssd1 vccd1 vccd1 _2850_/S sky130_fd_sc_hd__clkbuf_2
X_2767_ _2767_/A _2767_/B vssd1 vssd1 vccd1 vccd1 _2768_/A sky130_fd_sc_hd__and2_1
X_2698_ _2982_/A vssd1 vssd1 vccd1 vccd1 _2769_/A sky130_fd_sc_hd__buf_2
X_4506_ _4506_/A vssd1 vssd1 vccd1 vccd1 _5056_/D sky130_fd_sc_hd__clkbuf_1
X_4437_ _4454_/A vssd1 vssd1 vccd1 vccd1 _4452_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _5022_/Q _4315_/X _4367_/Y _2869_/X vssd1 vssd1 vccd1 vccd1 _5022_/D sky130_fd_sc_hd__o211a_1
X_3319_ _3327_/A vssd1 vssd1 vccd1 vccd1 _3320_/A sky130_fd_sc_hd__clkinv_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4290_/A _4292_/Y _4297_/X _4230_/A vssd1 vssd1 vccd1 vccd1 _4299_/X sky130_fd_sc_hd__a31o_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3670_ _5114_/Q _4946_/Q vssd1 vssd1 vccd1 vccd1 _3671_/B sky130_fd_sc_hd__or2_1
X_2621_ _2621_/A vssd1 vssd1 vccd1 vccd1 _4753_/D sky130_fd_sc_hd__clkbuf_1
X_2552_ _3168_/A vssd1 vssd1 vccd1 vccd1 _4632_/A sky130_fd_sc_hd__clkbuf_4
X_5271_ _5271_/A _2464_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
X_2483_ _2484_/A vssd1 vssd1 vccd1 vccd1 _2483_/Y sky130_fd_sc_hd__inv_2
X_4222_ _5016_/Q _4796_/Q vssd1 vssd1 vccd1 vccd1 _4229_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4153_ _4144_/A _4146_/Y _4151_/Y _4136_/X vssd1 vssd1 vccd1 vccd1 _4153_/X sky130_fd_sc_hd__a31o_1
X_4084_ _4998_/Q _4778_/Q vssd1 vssd1 vccd1 vccd1 _4084_/Y sky130_fd_sc_hd__nand2_1
X_3104_ _4876_/Q _5044_/Q vssd1 vssd1 vccd1 vccd1 _3105_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3035_ _3032_/Y _3026_/X _3039_/B _3041_/C vssd1 vssd1 vccd1 vccd1 _3035_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4986_ _4989_/CLK _4986_/D vssd1 vssd1 vccd1 vccd1 _4986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3937_ _3943_/A vssd1 vssd1 vccd1 vccd1 _3937_/X sky130_fd_sc_hd__buf_2
X_3868_ _4972_/Q _4752_/Q vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__and2_1
X_2819_ _4441_/A vssd1 vssd1 vccd1 vccd1 _2833_/S sky130_fd_sc_hd__clkbuf_2
X_3799_ _4963_/Q _4743_/Q vssd1 vssd1 vccd1 vccd1 _3805_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5199__106 vssd1 vssd1 vccd1 vccd1 _5199__106/HI _5307_/A sky130_fd_sc_hd__conb_1
XFILLER_74_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 la1_data_in[20] vssd1 vssd1 vccd1 vccd1 _2858_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput29 la1_data_in[31] vssd1 vssd1 vccd1 vccd1 _2905_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4840_ _5041_/CLK _4840_/D vssd1 vssd1 vccd1 vccd1 _5281_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _5018_/CLK _4771_/D vssd1 vssd1 vccd1 vccd1 _4771_/Q sky130_fd_sc_hd__dfxtp_1
X_3722_ _3722_/A _3722_/B vssd1 vssd1 vccd1 vccd1 _3722_/Y sky130_fd_sc_hd__nand2_2
X_3653_ _5112_/Q _4944_/Q vssd1 vssd1 vccd1 vccd1 _3663_/A sky130_fd_sc_hd__nand2_1
X_2604_ _4957_/Q _4749_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _2605_/B sky130_fd_sc_hd__mux2_1
X_5323_ _5323_/A _2526_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
X_3584_ _4936_/Q _5104_/Q vssd1 vssd1 vccd1 vccd1 _3586_/A sky130_fd_sc_hd__and2_1
X_2535_ _2539_/A vssd1 vssd1 vccd1 vccd1 _2535_/Y sky130_fd_sc_hd__inv_2
X_2466_ _2466_/A vssd1 vssd1 vccd1 vccd1 _2466_/Y sky130_fd_sc_hd__inv_2
X_5254_ _5254_/A _2443_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
X_4205_ _4196_/A _4198_/Y _4203_/X _4136_/A vssd1 vssd1 vccd1 vccd1 _4205_/X sky130_fd_sc_hd__a31o_1
X_4136_ _4136_/A vssd1 vssd1 vccd1 vccd1 _4136_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ _4093_/A _4067_/B vssd1 vssd1 vccd1 vccd1 _4067_/X sky130_fd_sc_hd__xor2_1
XFILLER_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3018_ _4865_/Q _5033_/Q vssd1 vssd1 vccd1 vccd1 _3019_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4969_ _4972_/CLK _4969_/D vssd1 vssd1 vccd1 vccd1 _4969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4836_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4823_ _5050_/CLK _4823_/D vssd1 vssd1 vccd1 vccd1 _4823_/Q sky130_fd_sc_hd__dfxtp_1
X_4754_ _4966_/CLK _4754_/D vssd1 vssd1 vccd1 vccd1 _4754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ _5119_/Q _4951_/Q vssd1 vssd1 vccd1 vccd1 _3711_/B sky130_fd_sc_hd__nand2_1
X_4685_ _4702_/A vssd1 vssd1 vccd1 vccd1 _4699_/S sky130_fd_sc_hd__buf_2
X_3636_ _3636_/A _3636_/B vssd1 vssd1 vccd1 vccd1 _3638_/A sky130_fd_sc_hd__or2_1
X_3567_ _4921_/Q _3554_/X _3565_/X _3566_/X vssd1 vssd1 vccd1 vccd1 _4921_/D sky130_fd_sc_hd__o211a_1
X_5306_ _5306_/A _2506_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
X_2518_ _2521_/A vssd1 vssd1 vccd1 vccd1 _2518_/Y sky130_fd_sc_hd__inv_2
X_3498_ _4925_/Q _5093_/Q vssd1 vssd1 vccd1 vccd1 _3500_/A sky130_fd_sc_hd__nor2_1
X_5237_ _5237_/A _2532_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2449_ _2453_/A vssd1 vssd1 vccd1 vccd1 _2449_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5099_ _5099_/CLK _5099_/D vssd1 vssd1 vccd1 vccd1 _5099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4119_ _4991_/Q vssd1 vssd1 vccd1 vccd1 _4119_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4470_ _4470_/A _4470_/B vssd1 vssd1 vccd1 vccd1 _4471_/A sky130_fd_sc_hd__and2_1
X_3421_ _3421_/A _3421_/B _3421_/C vssd1 vssd1 vccd1 vccd1 _3422_/C sky130_fd_sc_hd__and3_1
X_3352_ _4894_/Q _3352_/B vssd1 vssd1 vccd1 vccd1 _3352_/X sky130_fd_sc_hd__or2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _4898_/Q _5066_/Q vssd1 vssd1 vccd1 vccd1 _3285_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5026_/CLK _5022_/D vssd1 vssd1 vccd1 vccd1 _5022_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4806_ _5015_/CLK _4806_/D vssd1 vssd1 vccd1 vccd1 _4806_/Q sky130_fd_sc_hd__dfxtp_1
X_2998_ _2998_/A _2998_/B vssd1 vssd1 vccd1 vccd1 _2998_/Y sky130_fd_sc_hd__nand2_1
X_4737_ _5114_/CLK _4737_/D vssd1 vssd1 vccd1 vccd1 _4737_/Q sky130_fd_sc_hd__dfxtp_1
X_4668_ _4702_/A vssd1 vssd1 vccd1 vccd1 _4682_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_79_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3619_ _4939_/Q _5107_/Q _3606_/Y _3617_/C _3618_/X vssd1 vssd1 vccd1 vccd1 _3619_/X
+ sky130_fd_sc_hd__a221o_1
X_4599_ _4903_/Q _5083_/Q _4612_/S vssd1 vssd1 vccd1 vccd1 _4600_/B sky130_fd_sc_hd__mux2_1
XFILLER_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3970_ _3971_/A _3971_/B vssd1 vssd1 vccd1 vccd1 _3970_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2921_ _2934_/A _2921_/B vssd1 vssd1 vccd1 vccd1 _2922_/A sky130_fd_sc_hd__and2_1
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2852_ _2852_/A vssd1 vssd1 vccd1 vccd1 _4819_/D sky130_fd_sc_hd__clkbuf_1
X_2783_ _5008_/Q _4800_/Q _2798_/S vssd1 vssd1 vccd1 vccd1 _2784_/B sky130_fd_sc_hd__mux2_1
X_4522_ _4522_/A _4522_/B vssd1 vssd1 vccd1 vccd1 _4523_/A sky130_fd_sc_hd__and2_1
X_4453_ _4453_/A vssd1 vssd1 vccd1 vccd1 _5041_/D sky130_fd_sc_hd__clkbuf_1
X_3404_ _4913_/Q _5081_/Q vssd1 vssd1 vccd1 vccd1 _3405_/B sky130_fd_sc_hd__nand2_1
X_4384_ _4384_/A _4384_/B vssd1 vssd1 vccd1 vccd1 _4386_/B sky130_fd_sc_hd__and2_1
X_3335_ _4904_/Q _5072_/Q vssd1 vssd1 vccd1 vccd1 _3336_/B sky130_fd_sc_hd__or2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _4032_/A _3553_/B vssd1 vssd1 vccd1 vccd1 _3352_/B sky130_fd_sc_hd__nor2_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5026_/CLK _5005_/D vssd1 vssd1 vccd1 vccd1 _5005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3197_ _3197_/A _3197_/B vssd1 vssd1 vccd1 vccd1 _3197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3120_ _3137_/A vssd1 vssd1 vccd1 vccd1 _3120_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3051_ _4869_/Q _5037_/Q vssd1 vssd1 vccd1 vccd1 _3051_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3953_ _3954_/A _3954_/B vssd1 vssd1 vccd1 vccd1 _3953_/X sky130_fd_sc_hd__or2_1
XFILLER_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3884_ _3883_/A _3902_/B _3848_/X vssd1 vssd1 vccd1 vccd1 _3884_/X sky130_fd_sc_hd__a21o_1
X_2904_ _2855_/A _4830_/Q _2902_/X _2903_/X _2897_/X vssd1 vssd1 vccd1 vccd1 _4830_/D
+ sky130_fd_sc_hd__o221a_1
X_2835_ _2835_/A vssd1 vssd1 vccd1 vccd1 _4814_/D sky130_fd_sc_hd__clkbuf_1
X_2766_ _5003_/Q _4795_/Q _2779_/S vssd1 vssd1 vccd1 vccd1 _2767_/B sky130_fd_sc_hd__mux2_1
X_2697_ _2697_/A vssd1 vssd1 vccd1 vccd1 _4775_/D sky130_fd_sc_hd__clkbuf_1
X_4505_ _4505_/A _4505_/B vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__and2_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4436_ _4436_/A vssd1 vssd1 vccd1 vccd1 _5036_/D sky130_fd_sc_hd__clkbuf_1
X_4367_ _4367_/A _4367_/B vssd1 vssd1 vccd1 vccd1 _4367_/Y sky130_fd_sc_hd__nand2_1
X_3318_ _4902_/Q _5070_/Q vssd1 vssd1 vccd1 vccd1 _3318_/Y sky130_fd_sc_hd__nand2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4290_/A _4292_/Y _4297_/X vssd1 vssd1 vccd1 vccd1 _4298_/Y sky130_fd_sc_hd__a21oi_1
X_3249_ _3241_/A _3245_/X _3248_/X vssd1 vssd1 vccd1 vccd1 _3249_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5201__108 vssd1 vssd1 vccd1 vccd1 _5201__108/HI _5309_/A sky130_fd_sc_hd__conb_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ _2627_/A _2620_/B vssd1 vssd1 vccd1 vccd1 _2621_/A sky130_fd_sc_hd__and2_1
X_2551_ _2982_/A vssd1 vssd1 vccd1 vccd1 _2557_/A sky130_fd_sc_hd__buf_2
X_5270_ _5270_/A _2463_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
X_2482_ _2484_/A vssd1 vssd1 vccd1 vccd1 _2482_/Y sky130_fd_sc_hd__inv_2
X_4221_ _5016_/Q _4796_/Q vssd1 vssd1 vccd1 vccd1 _4221_/X sky130_fd_sc_hd__or2_1
X_4152_ _4144_/A _4146_/Y _4151_/Y vssd1 vssd1 vccd1 vccd1 _4152_/Y sky130_fd_sc_hd__a21oi_1
X_4083_ _4038_/X _4080_/Y _4081_/X _4082_/X vssd1 vssd1 vccd1 vccd1 _4986_/D sky130_fd_sc_hd__o211a_1
X_3103_ _4876_/Q _5044_/Q vssd1 vssd1 vccd1 vccd1 _3105_/A sky130_fd_sc_hd__and2_1
X_3034_ _4867_/Q _5035_/Q vssd1 vssd1 vccd1 vccd1 _3041_/C sky130_fd_sc_hd__or2_1
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4985_ _4989_/CLK _4985_/D vssd1 vssd1 vccd1 vccd1 _4985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3936_ _3936_/A _3936_/B vssd1 vssd1 vccd1 vccd1 _3943_/A sky130_fd_sc_hd__or2_2
X_3867_ _4959_/Q _3838_/X _3864_/Y _3865_/X _3866_/X vssd1 vssd1 vccd1 vccd1 _4959_/D
+ sky130_fd_sc_hd__o221a_1
X_2818_ _4632_/A vssd1 vssd1 vccd1 vccd1 _4441_/A sky130_fd_sc_hd__buf_2
X_3798_ _4950_/Q _3745_/X _3796_/X _3797_/X vssd1 vssd1 vccd1 vccd1 _4950_/D sky130_fd_sc_hd__o211a_1
X_2749_ _4998_/Q _4790_/Q _2762_/S vssd1 vssd1 vccd1 vccd1 _2750_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4419_ _4419_/A vssd1 vssd1 vccd1 vccd1 _5031_/D sky130_fd_sc_hd__clkbuf_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5114_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput19 la1_data_in[21] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4770_ _5018_/CLK _4770_/D vssd1 vssd1 vccd1 vccd1 _4770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ _3722_/A _3722_/B vssd1 vssd1 vccd1 vccd1 _3721_/X sky130_fd_sc_hd__or2_1
X_3652_ _3737_/B vssd1 vssd1 vccd1 vccd1 _3652_/X sky130_fd_sc_hd__clkbuf_2
X_2603_ _2603_/A vssd1 vssd1 vccd1 vccd1 _4748_/D sky130_fd_sc_hd__clkbuf_1
X_3583_ _4923_/Q _3554_/X _3581_/Y _3582_/X _3551_/X vssd1 vssd1 vccd1 vccd1 _4923_/D
+ sky130_fd_sc_hd__o221a_1
X_5322_ _5322_/A _2525_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
X_2534_ _2540_/A vssd1 vssd1 vccd1 vccd1 _2539_/A sky130_fd_sc_hd__buf_8
X_5253_ _5253_/A _2441_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
X_2465_ _2466_/A vssd1 vssd1 vccd1 vccd1 _2465_/Y sky130_fd_sc_hd__inv_2
X_4204_ _4196_/A _4198_/Y _4203_/X vssd1 vssd1 vccd1 vccd1 _4204_/Y sky130_fd_sc_hd__a21oi_1
X_4135_ _4135_/A _4135_/B vssd1 vssd1 vccd1 vccd1 _4135_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ _4051_/A _4051_/B _4057_/Y _4065_/X vssd1 vssd1 vccd1 vccd1 _4067_/B sky130_fd_sc_hd__a31o_1
X_3017_ _4865_/Q _5033_/Q vssd1 vssd1 vccd1 vccd1 _3019_/A sky130_fd_sc_hd__or2_1
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4968_ _4972_/CLK _4968_/D vssd1 vssd1 vccd1 vccd1 _4968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4899_ _5079_/CLK _4899_/D vssd1 vssd1 vccd1 vccd1 _4899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3919_ _4978_/Q _4758_/Q vssd1 vssd1 vccd1 vccd1 _3921_/A sky130_fd_sc_hd__nor2_1
X_5207__114 vssd1 vssd1 vccd1 vccd1 _5207__114/HI _5315_/A sky130_fd_sc_hd__conb_1
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4822_ _5019_/CLK _4822_/D vssd1 vssd1 vccd1 vccd1 _4822_/Q sky130_fd_sc_hd__dfxtp_1
X_4753_ _4966_/CLK _4753_/D vssd1 vssd1 vccd1 vccd1 _4753_/Q sky130_fd_sc_hd__dfxtp_1
X_5169__76 vssd1 vssd1 vccd1 vccd1 _5169__76/HI _5264_/A sky130_fd_sc_hd__conb_1
X_3704_ _4938_/Q _3652_/X _3703_/X _3659_/X vssd1 vssd1 vccd1 vccd1 _4938_/D sky130_fd_sc_hd__o211a_1
X_4684_ _4684_/A vssd1 vssd1 vccd1 vccd1 _5107_/D sky130_fd_sc_hd__clkbuf_1
X_3635_ _4942_/Q _5110_/Q vssd1 vssd1 vccd1 vccd1 _3636_/B sky130_fd_sc_hd__and2_1
X_3566_ _3566_/A vssd1 vssd1 vccd1 vccd1 _3566_/X sky130_fd_sc_hd__clkbuf_2
X_2517_ _2521_/A vssd1 vssd1 vccd1 vccd1 _2517_/Y sky130_fd_sc_hd__inv_2
X_5305_ _5305_/A _2505_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_3497_ _3494_/A _3494_/B _3489_/A vssd1 vssd1 vccd1 vccd1 _3501_/A sky130_fd_sc_hd__a21oi_1
X_5236_ _5236_/A _2531_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
X_2448_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2453_/A sky130_fd_sc_hd__buf_8
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5098_ _5098_/CLK _5098_/D vssd1 vssd1 vccd1 vccd1 _5098_/Q sky130_fd_sc_hd__dfxtp_1
X_4118_ _4038_/X _4116_/X _4117_/X _4082_/X vssd1 vssd1 vccd1 vccd1 _4990_/D sky130_fd_sc_hd__o211a_1
X_4049_ _4049_/A _4049_/B vssd1 vssd1 vccd1 vccd1 _4051_/B sky130_fd_sc_hd__and2_1
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5183__90 vssd1 vssd1 vccd1 vccd1 _5183__90/HI _5291_/A sky130_fd_sc_hd__conb_1
XFILLER_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3420_ _4903_/Q _3401_/X _3418_/Y _3419_/X _3325_/X vssd1 vssd1 vccd1 vccd1 _4903_/D
+ sky130_fd_sc_hd__o221a_1
X_3351_ _3351_/A _3351_/B vssd1 vssd1 vccd1 vccd1 _3351_/X sky130_fd_sc_hd__xor2_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3276_/A _3276_/B _3281_/Y vssd1 vssd1 vccd1 vccd1 _3287_/A sky130_fd_sc_hd__o21ai_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5021_ _5026_/CLK _5021_/D vssd1 vssd1 vccd1 vccd1 _5021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4805_ _5015_/CLK _4805_/D vssd1 vssd1 vccd1 vccd1 _4805_/Q sky130_fd_sc_hd__dfxtp_1
X_2997_ _2998_/A _2998_/B vssd1 vssd1 vccd1 vccd1 _2997_/X sky130_fd_sc_hd__or2_1
X_4736_ _5114_/CLK _4736_/D vssd1 vssd1 vccd1 vccd1 _4736_/Q sky130_fd_sc_hd__dfxtp_1
X_4667_ _4667_/A vssd1 vssd1 vccd1 vccd1 _5102_/D sky130_fd_sc_hd__clkbuf_1
X_3618_ _4938_/Q _5106_/Q _3618_/C vssd1 vssd1 vccd1 vccd1 _3618_/X sky130_fd_sc_hd__and3_1
X_4598_ _4615_/A vssd1 vssd1 vccd1 vccd1 _4612_/S sky130_fd_sc_hd__clkbuf_2
X_3549_ _3541_/B _3547_/X _3548_/X vssd1 vssd1 vccd1 vccd1 _3549_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5219_ _5219_/A _2419_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_29_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2920_ _5274_/A _4849_/Q _2968_/B vssd1 vssd1 vccd1 vccd1 _2921_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2851_ _2917_/A _2851_/B vssd1 vssd1 vccd1 vccd1 _2852_/A sky130_fd_sc_hd__and2_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2782_ _2801_/A vssd1 vssd1 vccd1 vccd1 _2798_/S sky130_fd_sc_hd__clkbuf_2
X_4521_ _4881_/Q _5061_/Q _4525_/S vssd1 vssd1 vccd1 vccd1 _4522_/B sky130_fd_sc_hd__mux2_1
X_5139__46 vssd1 vssd1 vccd1 vccd1 _5139__46/HI _5234_/A sky130_fd_sc_hd__conb_1
X_4452_ _4452_/A _4452_/B vssd1 vssd1 vccd1 vccd1 _4453_/A sky130_fd_sc_hd__and2_1
X_3403_ _4913_/Q _5081_/Q vssd1 vssd1 vccd1 vccd1 _3403_/Y sky130_fd_sc_hd__nor2_1
X_4383_ _4828_/Q _4816_/Q vssd1 vssd1 vccd1 vccd1 _4384_/B sky130_fd_sc_hd__or2_1
X_3334_ _4904_/Q _5072_/Q vssd1 vssd1 vccd1 vccd1 _3336_/A sky130_fd_sc_hd__nand2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3265_ _3557_/B vssd1 vssd1 vccd1 vccd1 _3553_/B sky130_fd_sc_hd__clkbuf_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5004_/CLK _5004_/D vssd1 vssd1 vccd1 vccd1 _5004_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _4887_/Q _5055_/Q vssd1 vssd1 vccd1 vccd1 _3197_/B sky130_fd_sc_hd__and2_1
XFILLER_81_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4719_ _4719_/A vssd1 vssd1 vccd1 vccd1 _4732_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5041_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5153__60 vssd1 vssd1 vccd1 vccd1 _5153__60/HI _5248_/A sky130_fd_sc_hd__conb_1
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3050_ _4856_/Q _2976_/X _3049_/X _2983_/X vssd1 vssd1 vccd1 vccd1 _4856_/D sky130_fd_sc_hd__o211a_1
XFILLER_63_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3952_ _3952_/A _3952_/B vssd1 vssd1 vccd1 vccd1 _3954_/B sky130_fd_sc_hd__and2_1
X_3883_ _3883_/A _3902_/B vssd1 vssd1 vccd1 vccd1 _3883_/Y sky130_fd_sc_hd__nor2_1
X_2903_ _2889_/X input28/X _2958_/B vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__a21bo_1
X_2834_ _2838_/A _2834_/B vssd1 vssd1 vccd1 vccd1 _2835_/A sky130_fd_sc_hd__and2_1
X_2765_ _2801_/A vssd1 vssd1 vccd1 vccd1 _2779_/S sky130_fd_sc_hd__buf_2
X_4504_ _4876_/Q _5056_/Q _4508_/S vssd1 vssd1 vccd1 vccd1 _4505_/B sky130_fd_sc_hd__mux2_1
X_2696_ _2696_/A _2696_/B vssd1 vssd1 vccd1 vccd1 _2697_/A sky130_fd_sc_hd__and2_1
X_4435_ _4435_/A _4435_/B vssd1 vssd1 vccd1 vccd1 _4436_/A sky130_fd_sc_hd__and2_1
X_4366_ _4369_/A _4369_/B vssd1 vssd1 vccd1 vccd1 _4367_/B sky130_fd_sc_hd__xnor2_1
X_3317_ _3272_/X _3315_/Y _3316_/X _3279_/X vssd1 vssd1 vccd1 vccd1 _4890_/D sky130_fd_sc_hd__o211a_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4295_/Y _4297_/B vssd1 vssd1 vccd1 vccd1 _4297_/X sky130_fd_sc_hd__and2b_1
XFILLER_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3248_ _3246_/Y _3248_/B vssd1 vssd1 vccd1 vccd1 _3248_/X sky130_fd_sc_hd__and2b_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3179_ _4885_/Q _5053_/Q vssd1 vssd1 vccd1 vccd1 _3181_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ _3133_/A vssd1 vssd1 vccd1 vccd1 _2982_/A sky130_fd_sc_hd__clkbuf_2
X_2481_ _2484_/A vssd1 vssd1 vccd1 vccd1 _2481_/Y sky130_fd_sc_hd__inv_2
X_4220_ _4306_/B vssd1 vssd1 vccd1 vccd1 _4220_/X sky130_fd_sc_hd__clkbuf_2
X_4151_ _4151_/A _4151_/B vssd1 vssd1 vccd1 vccd1 _4151_/Y sky130_fd_sc_hd__nor2_1
X_3102_ _4863_/Q _3074_/X _3100_/Y _3101_/X _3037_/X vssd1 vssd1 vccd1 vccd1 _4863_/D
+ sky130_fd_sc_hd__o221a_1
X_4082_ _4321_/A vssd1 vssd1 vccd1 vccd1 _4082_/X sky130_fd_sc_hd__clkbuf_2
X_3033_ _4867_/Q _5035_/Q vssd1 vssd1 vccd1 vccd1 _3039_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4984_ _4989_/CLK _4984_/D vssd1 vssd1 vccd1 vccd1 _4984_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3935_ _4980_/Q _4760_/Q vssd1 vssd1 vccd1 vccd1 _3942_/A sky130_fd_sc_hd__nand2_1
X_3866_ _4076_/A vssd1 vssd1 vccd1 vccd1 _3866_/X sky130_fd_sc_hd__clkbuf_2
X_3797_ _3945_/A vssd1 vssd1 vccd1 vccd1 _3797_/X sky130_fd_sc_hd__buf_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2817_ _2817_/A vssd1 vssd1 vccd1 vccd1 _4809_/D sky130_fd_sc_hd__clkbuf_1
X_2748_ _2801_/A vssd1 vssd1 vccd1 vccd1 _2762_/S sky130_fd_sc_hd__clkbuf_2
X_4418_ _4418_/A _4418_/B vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__and2_1
X_2679_ _2679_/A _2679_/B vssd1 vssd1 vccd1 vccd1 _2680_/A sky130_fd_sc_hd__and2_1
X_5123__30 vssd1 vssd1 vccd1 vccd1 _5123__30/HI _5218_/A sky130_fd_sc_hd__conb_1
X_4349_ _4822_/Q _4810_/Q _4348_/X _4341_/B vssd1 vssd1 vccd1 vccd1 _4349_/X sky130_fd_sc_hd__a31o_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3720_ _3720_/A _3720_/B vssd1 vssd1 vccd1 vccd1 _3722_/B sky130_fd_sc_hd__and2_1
XFILLER_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3651_ _3651_/A vssd1 vssd1 vccd1 vccd1 _3737_/B sky130_fd_sc_hd__clkbuf_2
X_2602_ _2609_/A _2602_/B vssd1 vssd1 vccd1 vccd1 _2603_/A sky130_fd_sc_hd__and2_1
X_3582_ _3573_/A _3575_/Y _3580_/Y _3564_/X vssd1 vssd1 vccd1 vccd1 _3582_/X sky130_fd_sc_hd__a31o_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5321_ _5321_/A _2524_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
X_2533_ _2533_/A vssd1 vssd1 vccd1 vccd1 _2533_/Y sky130_fd_sc_hd__inv_2
X_2464_ _2466_/A vssd1 vssd1 vccd1 vccd1 _2464_/Y sky130_fd_sc_hd__inv_2
X_5252_ _5252_/A _2440_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
X_4203_ _4201_/Y _4203_/B vssd1 vssd1 vccd1 vccd1 _4203_/X sky130_fd_sc_hd__and2b_1
X_4134_ _4135_/A _4135_/B vssd1 vssd1 vccd1 vccd1 _4134_/X sky130_fd_sc_hd__or2_1
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4065_ _4994_/Q _4774_/Q _4064_/X _4057_/B vssd1 vssd1 vccd1 vccd1 _4065_/X sky130_fd_sc_hd__a31o_1
X_3016_ _3040_/A _3013_/B _3009_/A vssd1 vssd1 vccd1 vccd1 _3020_/A sky130_fd_sc_hd__a21oi_1
XFILLER_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _4978_/CLK _4967_/D vssd1 vssd1 vccd1 vccd1 _4967_/Q sky130_fd_sc_hd__dfxtp_1
X_3918_ _4965_/Q _3878_/X _3916_/Y _3917_/X _3866_/X vssd1 vssd1 vccd1 vccd1 _4965_/D
+ sky130_fd_sc_hd__o221a_1
X_4898_ _5077_/CLK _4898_/D vssd1 vssd1 vccd1 vccd1 _4898_/Q sky130_fd_sc_hd__dfxtp_1
X_3849_ _3846_/X _3847_/Y _3848_/X vssd1 vssd1 vccd1 vccd1 _3849_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4821_ _5019_/CLK _4821_/D vssd1 vssd1 vccd1 vccd1 _4821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4752_ _4752_/CLK _4752_/D vssd1 vssd1 vccd1 vccd1 _4752_/Q sky130_fd_sc_hd__dfxtp_1
X_4683_ _4696_/A _4683_/B vssd1 vssd1 vccd1 vccd1 _4684_/A sky130_fd_sc_hd__and2_1
X_3703_ _3701_/Y _3702_/X _3680_/X vssd1 vssd1 vccd1 vccd1 _3703_/X sky130_fd_sc_hd__a21o_1
X_3634_ _4942_/Q _5110_/Q vssd1 vssd1 vccd1 vccd1 _3636_/A sky130_fd_sc_hd__nor2_1
X_3565_ _3562_/X _3563_/Y _3564_/X vssd1 vssd1 vccd1 vccd1 _3565_/X sky130_fd_sc_hd__a21o_1
X_2516_ _2516_/A vssd1 vssd1 vccd1 vccd1 _2521_/A sky130_fd_sc_hd__buf_8
X_5304_ _5304_/A _2503_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
X_3496_ _4912_/Q _3457_/X _3495_/X _3434_/X vssd1 vssd1 vccd1 vccd1 _4912_/D sky130_fd_sc_hd__o211a_1
X_5235_ _5235_/A _2530_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
X_2447_ _2447_/A vssd1 vssd1 vccd1 vccd1 _2447_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5097_ _5107_/CLK _5097_/D vssd1 vssd1 vccd1 vccd1 _5097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4117_ _4990_/Q _4117_/B vssd1 vssd1 vccd1 vccd1 _4117_/X sky130_fd_sc_hd__or2_1
X_4048_ _4994_/Q _4774_/Q vssd1 vssd1 vccd1 vccd1 _4049_/B sky130_fd_sc_hd__or2_1
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3350_ _3336_/A _3338_/Y _3343_/B _3341_/Y vssd1 vssd1 vccd1 vccd1 _3351_/B sky130_fd_sc_hd__a31o_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _4897_/Q _5065_/Q vssd1 vssd1 vccd1 vccd1 _3281_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5020_ _5026_/CLK _5020_/D vssd1 vssd1 vccd1 vccd1 _5020_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4804_ _5015_/CLK _4804_/D vssd1 vssd1 vccd1 vccd1 _4804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2996_ _2996_/A _2996_/B vssd1 vssd1 vccd1 vccd1 _2998_/B sky130_fd_sc_hd__and2_1
X_4735_ _5122_/CLK _4735_/D vssd1 vssd1 vccd1 vccd1 _4735_/Q sky130_fd_sc_hd__dfxtp_1
X_4666_ _4679_/A _4666_/B vssd1 vssd1 vccd1 vccd1 _4667_/A sky130_fd_sc_hd__and2_1
X_4597_ _4597_/A vssd1 vssd1 vccd1 vccd1 _5082_/D sky130_fd_sc_hd__clkbuf_1
X_3617_ _3617_/A _3617_/B _3617_/C vssd1 vssd1 vccd1 vccd1 _3617_/X sky130_fd_sc_hd__and3_1
X_3548_ _4931_/Q _5099_/Q vssd1 vssd1 vccd1 vccd1 _3548_/X sky130_fd_sc_hd__xor2_1
X_3479_ _5285_/A vssd1 vssd1 vccd1 vccd1 _3479_/X sky130_fd_sc_hd__buf_2
X_5218_ _5218_/A _2418_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_28_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2850_ _5027_/Q _4819_/Q _2850_/S vssd1 vssd1 vccd1 vccd1 _2851_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2781_ _2781_/A vssd1 vssd1 vccd1 vccd1 _4799_/D sky130_fd_sc_hd__clkbuf_1
X_4520_ _4520_/A vssd1 vssd1 vccd1 vccd1 _5060_/D sky130_fd_sc_hd__clkbuf_1
X_4451_ _4861_/Q _5041_/Q _4455_/S vssd1 vssd1 vccd1 vccd1 _4452_/B sky130_fd_sc_hd__mux2_1
X_3402_ _3422_/A _3398_/B _3394_/A vssd1 vssd1 vccd1 vccd1 _3406_/A sky130_fd_sc_hd__a21oi_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4382_ _4828_/Q _4816_/Q vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__nand2_1
X_3333_ _3303_/B _3328_/X _3332_/X vssd1 vssd1 vccd1 vccd1 _3338_/A sky130_fd_sc_hd__a21o_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _4846_/Q _3648_/A vssd1 vssd1 vccd1 vccd1 _3557_/B sky130_fd_sc_hd__or2b_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5010_/CLK _5003_/D vssd1 vssd1 vccd1 vccd1 _5003_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _4887_/Q _5055_/Q vssd1 vssd1 vccd1 vccd1 _3197_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2979_ _3175_/A _4129_/A vssd1 vssd1 vccd1 vccd1 _2988_/A sky130_fd_sc_hd__or2_2
X_4718_ _4718_/A vssd1 vssd1 vccd1 vccd1 _5117_/D sky130_fd_sc_hd__clkbuf_1
X_4649_ _4662_/A _4649_/B vssd1 vssd1 vccd1 vccd1 _4650_/A sky130_fd_sc_hd__and2_1
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_18_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4981_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3951_ _4982_/Q _4762_/Q vssd1 vssd1 vccd1 vccd1 _3952_/B sky130_fd_sc_hd__or2_1
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2902_ _2886_/X input13/X _2887_/X vssd1 vssd1 vccd1 vccd1 _2902_/X sky130_fd_sc_hd__o21a_1
X_3882_ _3882_/A _3882_/B vssd1 vssd1 vccd1 vccd1 _3902_/B sky130_fd_sc_hd__and2_1
XFILLER_31_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2833_ _5022_/Q _4814_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _2834_/B sky130_fd_sc_hd__mux2_1
X_2764_ _2764_/A vssd1 vssd1 vccd1 vccd1 _4794_/D sky130_fd_sc_hd__clkbuf_1
X_4503_ _4503_/A vssd1 vssd1 vccd1 vccd1 _5055_/D sky130_fd_sc_hd__clkbuf_1
X_2695_ _4983_/Q _4775_/Q _2710_/S vssd1 vssd1 vccd1 vccd1 _2696_/B sky130_fd_sc_hd__mux2_1
X_4434_ _4856_/Q _5036_/Q _4438_/S vssd1 vssd1 vccd1 vccd1 _4435_/B sky130_fd_sc_hd__mux2_1
X_4365_ _4358_/A _4357_/B _4355_/Y vssd1 vssd1 vccd1 vccd1 _4369_/B sky130_fd_sc_hd__a21o_1
X_3316_ _4890_/Q _3352_/B vssd1 vssd1 vccd1 vccd1 _3316_/X sky130_fd_sc_hd__or2_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _5025_/Q _4805_/Q vssd1 vssd1 vccd1 vccd1 _4297_/B sky130_fd_sc_hd__nand2_1
X_3247_ _4893_/Q _5061_/Q vssd1 vssd1 vccd1 vccd1 _3248_/B sky130_fd_sc_hd__nand2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _4872_/Q _3172_/X _3177_/X _3148_/X vssd1 vssd1 vccd1 vccd1 _4872_/D sky130_fd_sc_hd__o211a_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2480_ _2484_/A vssd1 vssd1 vccd1 vccd1 _2480_/Y sky130_fd_sc_hd__inv_2
X_4150_ _5007_/Q _4787_/Q vssd1 vssd1 vccd1 vccd1 _4151_/B sky130_fd_sc_hd__and2_1
X_3101_ _3092_/A _3094_/Y _3099_/Y _3084_/X vssd1 vssd1 vccd1 vccd1 _3101_/X sky130_fd_sc_hd__a31o_1
X_4081_ _4986_/Q _4117_/B vssd1 vssd1 vccd1 vccd1 _4081_/X sky130_fd_sc_hd__or2_1
X_3032_ _4866_/Q _5034_/Q vssd1 vssd1 vccd1 vccd1 _3032_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4983_ _4983_/CLK _4983_/D vssd1 vssd1 vccd1 vccd1 _4983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3934_ _4980_/Q _4760_/Q vssd1 vssd1 vccd1 vccd1 _3934_/X sky130_fd_sc_hd__or2_1
X_3865_ _3856_/A _3858_/Y _3863_/Y _3848_/X vssd1 vssd1 vccd1 vccd1 _3865_/X sky130_fd_sc_hd__a31o_1
X_2816_ _2821_/A _2816_/B vssd1 vssd1 vccd1 vccd1 _2817_/A sky130_fd_sc_hd__and2_1
X_3796_ _3794_/Y _3795_/X _3755_/X vssd1 vssd1 vccd1 vccd1 _3796_/X sky130_fd_sc_hd__a21o_1
X_2747_ _2747_/A vssd1 vssd1 vccd1 vccd1 _4789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2678_ _4978_/Q _4770_/Q _2691_/S vssd1 vssd1 vccd1 vccd1 _2679_/B sky130_fd_sc_hd__mux2_1
X_4417_ _4851_/Q _5031_/Q _4421_/S vssd1 vssd1 vccd1 vccd1 _4418_/B sky130_fd_sc_hd__mux2_1
X_4348_ _4823_/Q _4811_/Q vssd1 vssd1 vccd1 vccd1 _4348_/X sky130_fd_sc_hd__or2_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4279_ _4276_/Y _4270_/X _4283_/B _4285_/C vssd1 vssd1 vccd1 vccd1 _4279_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5091_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3650_ _4032_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _3651_/A sky130_fd_sc_hd__nor2_1
X_2601_ _4956_/Q _4748_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _2602_/B sky130_fd_sc_hd__mux2_1
X_3581_ _3573_/A _3575_/Y _3580_/Y vssd1 vssd1 vccd1 vccd1 _3581_/Y sky130_fd_sc_hd__a21oi_1
X_5320_ _5320_/A _2523_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
X_2532_ _2533_/A vssd1 vssd1 vccd1 vccd1 _2532_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5251_ _5251_/A _2439_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2463_ _2466_/A vssd1 vssd1 vccd1 vccd1 _2463_/Y sky130_fd_sc_hd__inv_2
X_4202_ _5013_/Q _4793_/Q vssd1 vssd1 vccd1 vccd1 _4203_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4133_ _5005_/Q _4785_/Q vssd1 vssd1 vccd1 vccd1 _4135_/B sky130_fd_sc_hd__xnor2_1
X_4064_ _4995_/Q _4775_/Q vssd1 vssd1 vccd1 vccd1 _4064_/X sky130_fd_sc_hd__or2_1
X_3015_ _2980_/X _3013_/X _3014_/X _2983_/X vssd1 vssd1 vccd1 vccd1 _4852_/D sky130_fd_sc_hd__o211a_1
XFILLER_24_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4966_ _4966_/CLK _4966_/D vssd1 vssd1 vccd1 vccd1 _4966_/Q sky130_fd_sc_hd__dfxtp_1
X_3917_ _3908_/A _3910_/Y _3915_/X _3848_/A vssd1 vssd1 vccd1 vccd1 _3917_/X sky130_fd_sc_hd__a31o_1
X_4897_ _5077_/CLK _4897_/D vssd1 vssd1 vccd1 vccd1 _4897_/Q sky130_fd_sc_hd__dfxtp_1
X_3848_ _3848_/A vssd1 vssd1 vccd1 vccd1 _3848_/X sky130_fd_sc_hd__clkbuf_2
X_3779_ _4958_/Q _4738_/Q _3778_/X _3770_/B vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__a31o_1
XFILLER_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4820_ _5019_/CLK _4820_/D vssd1 vssd1 vccd1 vccd1 _4820_/Q sky130_fd_sc_hd__dfxtp_1
X_4751_ _4752_/CLK _4751_/D vssd1 vssd1 vccd1 vccd1 _4751_/Q sky130_fd_sc_hd__dfxtp_1
X_4682_ _3517_/A _5107_/Q _4682_/S vssd1 vssd1 vccd1 vccd1 _4683_/B sky130_fd_sc_hd__mux2_1
X_3702_ _3711_/A _3702_/B vssd1 vssd1 vccd1 vccd1 _3702_/X sky130_fd_sc_hd__or2_1
X_3633_ _4929_/Q _3593_/X _3631_/Y _3632_/X _3551_/X vssd1 vssd1 vccd1 vccd1 _4929_/D
+ sky130_fd_sc_hd__o221a_1
X_3564_ _3564_/A vssd1 vssd1 vccd1 vccd1 _3564_/X sky130_fd_sc_hd__clkbuf_2
X_5303_ _5303_/A _2502_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
X_2515_ _2515_/A vssd1 vssd1 vccd1 vccd1 _2515_/Y sky130_fd_sc_hd__inv_2
X_3495_ _3493_/Y _3494_/X _3467_/X vssd1 vssd1 vccd1 vccd1 _3495_/X sky130_fd_sc_hd__a21o_1
X_5234_ _5234_/A _2438_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
X_2446_ _2447_/A vssd1 vssd1 vccd1 vccd1 _2446_/Y sky130_fd_sc_hd__inv_2
X_4116_ _4116_/A _4116_/B vssd1 vssd1 vccd1 vccd1 _4116_/X sky130_fd_sc_hd__xor2_1
X_5096_ _5107_/CLK _5096_/D vssd1 vssd1 vccd1 vccd1 _5096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4047_ _4994_/Q _4774_/Q vssd1 vssd1 vccd1 vccd1 _4049_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4949_ _4954_/CLK _4949_/D vssd1 vssd1 vccd1 vccd1 _4949_/Q sky130_fd_sc_hd__dfxtp_1
X_5213__120 vssd1 vssd1 vccd1 vccd1 _5213__120/HI _5321_/A sky130_fd_sc_hd__conb_1
XFILLER_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5174__81 vssd1 vssd1 vccd1 vccd1 _5174__81/HI _5269_/A sky130_fd_sc_hd__conb_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _4885_/Q _3268_/X _3277_/Y _3279_/X vssd1 vssd1 vccd1 vccd1 _4885_/D sky130_fd_sc_hd__o211a_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4803_ _5026_/CLK _4803_/D vssd1 vssd1 vccd1 vccd1 _4803_/Q sky130_fd_sc_hd__dfxtp_1
X_2995_ _4862_/Q _5030_/Q vssd1 vssd1 vccd1 vccd1 _2996_/B sky130_fd_sc_hd__or2_1
X_4734_ _4734_/A vssd1 vssd1 vccd1 vccd1 _5122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4665_ _4922_/Q _5102_/Q _4665_/S vssd1 vssd1 vccd1 vccd1 _4666_/B sky130_fd_sc_hd__mux2_1
X_4596_ _4609_/A _4596_/B vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__and2_1
X_3616_ _3616_/A _3616_/B _3618_/C vssd1 vssd1 vccd1 vccd1 _3617_/C sky130_fd_sc_hd__and3_1
X_3547_ _3528_/A _3530_/X _3535_/B _3546_/Y _3533_/Y vssd1 vssd1 vccd1 vccd1 _3547_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3478_ _3476_/X _3477_/Y _3461_/X vssd1 vssd1 vccd1 vccd1 _3478_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2429_ input1/X vssd1 vssd1 vccd1 vccd1 _2454_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _5079_/CLK _5079_/D vssd1 vssd1 vccd1 vccd1 _5079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2780_ _2784_/A _2780_/B vssd1 vssd1 vccd1 vccd1 _2781_/A sky130_fd_sc_hd__and2_1
XFILLER_7_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _4450_/A vssd1 vssd1 vccd1 vccd1 _5040_/D sky130_fd_sc_hd__clkbuf_1
X_3401_ _3448_/B vssd1 vssd1 vccd1 vccd1 _3401_/X sky130_fd_sc_hd__clkbuf_2
X_4381_ _4351_/B _4376_/X _4380_/X vssd1 vssd1 vccd1 vccd1 _4386_/A sky130_fd_sc_hd__a21o_1
X_3332_ _4903_/Q _5071_/Q _3330_/Y _3328_/C _3331_/X vssd1 vssd1 vccd1 vccd1 _3332_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _4883_/Q _3223_/A _3261_/Y _3262_/X _3230_/X vssd1 vssd1 vccd1 vccd1 _4883_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/CLK _5002_/D vssd1 vssd1 vccd1 vccd1 _5002_/Q sky130_fd_sc_hd__dfxtp_1
X_3194_ _3176_/X _3192_/X _3193_/X _3148_/X vssd1 vssd1 vccd1 vccd1 _4874_/D sky130_fd_sc_hd__o211a_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2978_ _4860_/Q _5028_/Q vssd1 vssd1 vccd1 vccd1 _2987_/A sky130_fd_sc_hd__nand2_1
X_4717_ _4730_/A _4717_/B vssd1 vssd1 vccd1 vccd1 _4718_/A sky130_fd_sc_hd__and2_1
X_4648_ _4917_/Q _5097_/Q _4648_/S vssd1 vssd1 vccd1 vccd1 _4649_/B sky130_fd_sc_hd__mux2_1
X_4579_ _4592_/A _4579_/B vssd1 vssd1 vccd1 vccd1 _4580_/A sky130_fd_sc_hd__and2_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5144__51 vssd1 vssd1 vccd1 vccd1 _5144__51/HI _5239_/A sky130_fd_sc_hd__conb_1
XFILLER_48_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3950_ _4982_/Q _4762_/Q vssd1 vssd1 vccd1 vccd1 _3952_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2901_ _2855_/A _4829_/Q _2899_/X _2900_/X _2897_/X vssd1 vssd1 vccd1 vccd1 _4829_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3881_ _4973_/Q _4753_/Q vssd1 vssd1 vccd1 vccd1 _3882_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2832_ _2832_/A vssd1 vssd1 vccd1 vccd1 _4813_/D sky130_fd_sc_hd__clkbuf_1
X_2763_ _2767_/A _2763_/B vssd1 vssd1 vccd1 vccd1 _2764_/A sky130_fd_sc_hd__and2_1
X_4502_ _4505_/A _4502_/B vssd1 vssd1 vccd1 vccd1 _4503_/A sky130_fd_sc_hd__and2_1
X_2694_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2710_/S sky130_fd_sc_hd__clkbuf_2
X_4433_ _4433_/A vssd1 vssd1 vccd1 vccd1 _5035_/D sky130_fd_sc_hd__clkbuf_1
X_4364_ _4375_/A _4375_/B vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__nand2_1
X_3315_ _3327_/A _3320_/B vssd1 vssd1 vccd1 vccd1 _3315_/Y sky130_fd_sc_hd__xnor2_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _5025_/Q _4805_/Q vssd1 vssd1 vccd1 vccd1 _4295_/Y sky130_fd_sc_hd__nor2_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _4893_/Q _5061_/Q vssd1 vssd1 vccd1 vccd1 _3246_/Y sky130_fd_sc_hd__nor2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3173_/X _3181_/A _3176_/X vssd1 vssd1 vccd1 vccd1 _3177_/X sky130_fd_sc_hd__a21o_1
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3100_ _3092_/A _3094_/Y _3099_/Y vssd1 vssd1 vccd1 vccd1 _3100_/Y sky130_fd_sc_hd__a21oi_1
X_4080_ _4092_/A _4086_/B vssd1 vssd1 vccd1 vccd1 _4080_/Y sky130_fd_sc_hd__xnor2_1
X_3031_ _4854_/Q _2976_/X _3030_/X _2983_/X vssd1 vssd1 vccd1 vccd1 _4854_/D sky130_fd_sc_hd__o211a_1
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4982_ _4983_/CLK _4982_/D vssd1 vssd1 vccd1 vccd1 _4982_/Q sky130_fd_sc_hd__dfxtp_1
X_3933_ _3933_/A vssd1 vssd1 vccd1 vccd1 _3933_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_3_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5019_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3864_ _3856_/A _3858_/Y _3863_/Y vssd1 vssd1 vccd1 vccd1 _3864_/Y sky130_fd_sc_hd__a21oi_1
X_2815_ _5017_/Q _4809_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _2816_/B sky130_fd_sc_hd__mux2_1
X_3795_ _3805_/A _3795_/B vssd1 vssd1 vccd1 vccd1 _3795_/X sky130_fd_sc_hd__or2_1
X_2746_ _2750_/A _2746_/B vssd1 vssd1 vccd1 vccd1 _2747_/A sky130_fd_sc_hd__and2_1
X_2677_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2691_/S sky130_fd_sc_hd__buf_2
X_4416_ _4416_/A vssd1 vssd1 vccd1 vccd1 _5030_/D sky130_fd_sc_hd__clkbuf_1
X_4347_ _4347_/A _4347_/B vssd1 vssd1 vccd1 vccd1 _4376_/A sky130_fd_sc_hd__nor2_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4278_ _5023_/Q _4803_/Q vssd1 vssd1 vccd1 vccd1 _4285_/C sky130_fd_sc_hd__or2_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _3232_/B _3225_/X _3232_/C _3236_/C _3182_/A vssd1 vssd1 vccd1 vccd1 _3229_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3580_ _3580_/A _3580_/B vssd1 vssd1 vccd1 vccd1 _3580_/Y sky130_fd_sc_hd__nor2_1
X_2600_ _2600_/A vssd1 vssd1 vccd1 vccd1 _4747_/D sky130_fd_sc_hd__clkbuf_1
X_2531_ _2533_/A vssd1 vssd1 vccd1 vccd1 _2531_/Y sky130_fd_sc_hd__inv_2
X_5250_ _5250_/A _2536_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_5_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4201_ _5013_/Q _4793_/Q vssd1 vssd1 vccd1 vccd1 _4201_/Y sky130_fd_sc_hd__nor2_1
X_2462_ _2466_/A vssd1 vssd1 vccd1 vccd1 _2462_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4132_ _4992_/Q _4126_/X _4131_/X _4082_/X vssd1 vssd1 vccd1 vccd1 _4992_/D sky130_fd_sc_hd__o211a_1
X_4063_ _4063_/A _4063_/B vssd1 vssd1 vccd1 vccd1 _4093_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3014_ _4852_/Q _3062_/B vssd1 vssd1 vccd1 vccd1 _3014_/X sky130_fd_sc_hd__or2_1
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4965_ _4966_/CLK _4965_/D vssd1 vssd1 vccd1 vccd1 _4965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3916_ _3908_/A _3910_/Y _3915_/X vssd1 vssd1 vccd1 vccd1 _3916_/Y sky130_fd_sc_hd__a21oi_1
X_4896_ _5077_/CLK _4896_/D vssd1 vssd1 vccd1 vccd1 _4896_/Q sky130_fd_sc_hd__dfxtp_1
X_3847_ _3847_/A _3847_/B vssd1 vssd1 vccd1 vccd1 _3847_/Y sky130_fd_sc_hd__nand2_1
X_3778_ _4959_/Q _4739_/Q vssd1 vssd1 vccd1 vccd1 _3778_/X sky130_fd_sc_hd__or2_1
X_2729_ _2729_/A vssd1 vssd1 vccd1 vccd1 _4784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4750_ _4964_/CLK _4750_/D vssd1 vssd1 vccd1 vccd1 _4750_/Q sky130_fd_sc_hd__dfxtp_1
X_4681_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4696_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3701_ _3711_/A _3702_/B vssd1 vssd1 vccd1 vccd1 _3701_/Y sky130_fd_sc_hd__nand2_1
X_3632_ _3623_/A _3625_/Y _3630_/X _3564_/A vssd1 vssd1 vccd1 vccd1 _3632_/X sky130_fd_sc_hd__a31o_1
X_5302_ _5302_/A _2501_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
X_3563_ _3563_/A _3563_/B vssd1 vssd1 vccd1 vccd1 _3563_/Y sky130_fd_sc_hd__nand2_1
X_2514_ _2515_/A vssd1 vssd1 vccd1 vccd1 _2514_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3494_ _3494_/A _3494_/B vssd1 vssd1 vccd1 vccd1 _3494_/X sky130_fd_sc_hd__or2_1
X_2445_ _2447_/A vssd1 vssd1 vccd1 vccd1 _2445_/Y sky130_fd_sc_hd__inv_2
X_5233_ _5233_/A _2437_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
X_4115_ _4101_/A _4103_/Y _4108_/B _4106_/Y vssd1 vssd1 vccd1 vccd1 _4116_/B sky130_fd_sc_hd__a31o_1
XFILLER_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5095_ _5107_/CLK _5095_/D vssd1 vssd1 vccd1 vccd1 _5095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4046_ _4042_/A _4042_/B _4045_/Y vssd1 vssd1 vccd1 vccd1 _4051_/A sky130_fd_sc_hd__o21ai_1
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4948_ _4948_/CLK _4948_/D vssd1 vssd1 vccd1 vccd1 _4948_/Q sky130_fd_sc_hd__dfxtp_1
X_4879_ _5087_/CLK _4879_/D vssd1 vssd1 vccd1 vccd1 _4879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5195__102 vssd1 vssd1 vccd1 vccd1 _5195__102/HI _5303_/A sky130_fd_sc_hd__conb_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2994_ _4862_/Q _5030_/Q vssd1 vssd1 vccd1 vccd1 _2996_/A sky130_fd_sc_hd__nand2_1
X_4802_ _5015_/CLK _4802_/D vssd1 vssd1 vccd1 vccd1 _4802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4733_ _4733_/A _4733_/B vssd1 vssd1 vccd1 vccd1 _4734_/A sky130_fd_sc_hd__and2_1
X_4664_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4679_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4595_ _4902_/Q _5082_/Q _4595_/S vssd1 vssd1 vccd1 vccd1 _4596_/B sky130_fd_sc_hd__mux2_1
X_3615_ _3517_/A _3593_/X _3613_/Y _3614_/X _3551_/X vssd1 vssd1 vccd1 vccd1 _4927_/D
+ sky130_fd_sc_hd__o221a_1
X_3546_ _3546_/A vssd1 vssd1 vccd1 vccd1 _3546_/Y sky130_fd_sc_hd__inv_2
X_3477_ _3477_/A _3477_/B vssd1 vssd1 vccd1 vccd1 _3477_/Y sky130_fd_sc_hd__nand2_1
X_2428_ _2428_/A vssd1 vssd1 vccd1 vccd1 _2428_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5078_ _5079_/CLK _5078_/D vssd1 vssd1 vccd1 vccd1 _5078_/Q sky130_fd_sc_hd__dfxtp_1
X_4029_ _4979_/Q _3933_/A _4027_/Y _4028_/X _3962_/X vssd1 vssd1 vccd1 vccd1 _4979_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3400_ _3367_/X _3398_/X _3399_/X _3353_/X vssd1 vssd1 vccd1 vccd1 _4900_/D sky130_fd_sc_hd__o211a_1
X_4380_ _4827_/Q _4815_/Q _4378_/Y _4376_/C _4379_/X vssd1 vssd1 vccd1 vccd1 _4380_/X
+ sky130_fd_sc_hd__a221o_1
X_3331_ _4902_/Q _5070_/Q _3331_/C vssd1 vssd1 vccd1 vccd1 _3331_/X sky130_fd_sc_hd__and3_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3254_/B _3259_/X _3260_/X _3182_/X vssd1 vssd1 vccd1 vccd1 _3262_/X sky130_fd_sc_hd__a31o_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5001_ _5010_/CLK _5001_/D vssd1 vssd1 vccd1 vccd1 _5001_/Q sky130_fd_sc_hd__dfxtp_1
X_3193_ _4874_/Q _3257_/B vssd1 vssd1 vccd1 vccd1 _3193_/X sky130_fd_sc_hd__or2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2977_ _4860_/Q _5028_/Q vssd1 vssd1 vccd1 vccd1 _2977_/X sky130_fd_sc_hd__or2_1
X_4716_ _4937_/Q _5117_/Q _4716_/S vssd1 vssd1 vccd1 vccd1 _4717_/B sky130_fd_sc_hd__mux2_1
X_4647_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4662_/A sky130_fd_sc_hd__clkbuf_2
X_4578_ _4897_/Q _5077_/Q _4578_/S vssd1 vssd1 vccd1 vccd1 _4579_/B sky130_fd_sc_hd__mux2_1
X_3529_ _3529_/A _3529_/B _3529_/C vssd1 vssd1 vccd1 vccd1 _3529_/Y sky130_fd_sc_hd__nand3_1
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5121_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2900_ _2889_/X input27/X _2883_/X vssd1 vssd1 vccd1 vccd1 _2900_/X sky130_fd_sc_hd__a21bo_1
X_3880_ _4973_/Q _4753_/Q vssd1 vssd1 vccd1 vccd1 _3882_/A sky130_fd_sc_hd__or2_1
XFILLER_31_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2831_ _2838_/A _2831_/B vssd1 vssd1 vccd1 vccd1 _2832_/A sky130_fd_sc_hd__and2_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2762_ _5002_/Q _4794_/Q _2762_/S vssd1 vssd1 vccd1 vccd1 _2763_/B sky130_fd_sc_hd__mux2_1
X_4501_ _4875_/Q _5055_/Q _4508_/S vssd1 vssd1 vccd1 vccd1 _4502_/B sky130_fd_sc_hd__mux2_1
X_2693_ _2693_/A vssd1 vssd1 vccd1 vccd1 _4774_/D sky130_fd_sc_hd__clkbuf_1
X_4432_ _4435_/A _4432_/B vssd1 vssd1 vccd1 vccd1 _4433_/A sky130_fd_sc_hd__and2_1
XANTENNA_0 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4363_ _4826_/Q _4814_/Q vssd1 vssd1 vccd1 vccd1 _4375_/B sky130_fd_sc_hd__nand2_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _3310_/A _3309_/B _3307_/Y vssd1 vssd1 vccd1 vccd1 _3320_/B sky130_fd_sc_hd__a21o_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _5012_/Q _4220_/X _4293_/X _4232_/X vssd1 vssd1 vccd1 vccd1 _5012_/D sky130_fd_sc_hd__o211a_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3245_/A _3242_/A vssd1 vssd1 vccd1 vccd1 _3245_/X sky130_fd_sc_hd__or2b_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3176_ _3182_/A vssd1 vssd1 vccd1 vccd1 _3176_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3030_ _3026_/X _3029_/X _2988_/X vssd1 vssd1 vccd1 vccd1 _3030_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _4981_/CLK _4981_/D vssd1 vssd1 vccd1 vccd1 _4981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3932_ _4021_/B vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__clkbuf_2
X_3863_ _3863_/A _3863_/B vssd1 vssd1 vccd1 vccd1 _3863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2814_ _2814_/A vssd1 vssd1 vccd1 vccd1 _4808_/D sky130_fd_sc_hd__clkbuf_1
X_3794_ _3805_/A _3795_/B vssd1 vssd1 vccd1 vccd1 _3794_/Y sky130_fd_sc_hd__nand2_1
X_2745_ _4997_/Q _4789_/Q _2745_/S vssd1 vssd1 vccd1 vccd1 _2746_/B sky130_fd_sc_hd__mux2_1
X_2676_ _2676_/A vssd1 vssd1 vccd1 vccd1 _4769_/D sky130_fd_sc_hd__clkbuf_1
X_4415_ _4418_/A _4415_/B vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__and2_1
X_4346_ _4824_/Q _4812_/Q vssd1 vssd1 vccd1 vccd1 _4347_/B sky130_fd_sc_hd__nor2_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4277_ _5023_/Q _4803_/Q vssd1 vssd1 vccd1 vccd1 _4283_/B sky130_fd_sc_hd__nand2_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ _3232_/B _3225_/X _3232_/C _3236_/C vssd1 vssd1 vccd1 vccd1 _3228_/Y sky130_fd_sc_hd__a22oi_1
X_3159_ _3144_/A _3146_/Y _3152_/B _3150_/Y vssd1 vssd1 vccd1 vccd1 _3160_/B sky130_fd_sc_hd__a31o_1
XFILLER_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_42_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5062_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2530_ _2533_/A vssd1 vssd1 vccd1 vccd1 _2530_/Y sky130_fd_sc_hd__inv_2
X_2461_ _2485_/A vssd1 vssd1 vccd1 vccd1 _2466_/A sky130_fd_sc_hd__buf_8
X_4200_ _5000_/Q _4126_/X _4199_/X _4163_/X vssd1 vssd1 vccd1 vccd1 _5000_/D sky130_fd_sc_hd__o211a_1
X_4131_ _4127_/X _4135_/A _4130_/X vssd1 vssd1 vccd1 vccd1 _4131_/X sky130_fd_sc_hd__a21o_1
X_4062_ _4996_/Q _4776_/Q vssd1 vssd1 vccd1 vccd1 _4063_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3013_ _3040_/A _3013_/B vssd1 vssd1 vccd1 vccd1 _3013_/X sky130_fd_sc_hd__xor2_1
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4964_ _4964_/CLK _4964_/D vssd1 vssd1 vccd1 vccd1 _4964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3915_ _3913_/Y _3915_/B vssd1 vssd1 vccd1 vccd1 _3915_/X sky130_fd_sc_hd__and2b_1
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4895_ _5099_/CLK _4895_/D vssd1 vssd1 vccd1 vccd1 _4895_/Q sky130_fd_sc_hd__dfxtp_1
X_3846_ _3847_/A _3847_/B vssd1 vssd1 vccd1 vccd1 _3846_/X sky130_fd_sc_hd__or2_1
X_3777_ _3777_/A _3777_/B vssd1 vssd1 vccd1 vccd1 _3806_/A sky130_fd_sc_hd__nor2_1
X_2728_ _2733_/A _2728_/B vssd1 vssd1 vccd1 vccd1 _2729_/A sky130_fd_sc_hd__and2_1
X_2659_ _2659_/A vssd1 vssd1 vccd1 vccd1 _4764_/D sky130_fd_sc_hd__clkbuf_1
X_4329_ _4821_/Q _4809_/Q vssd1 vssd1 vccd1 vccd1 _4329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3700_ _3692_/Y _3695_/B _3693_/Y vssd1 vssd1 vccd1 vccd1 _3702_/B sky130_fd_sc_hd__a21oi_1
X_4680_ _4680_/A vssd1 vssd1 vccd1 vccd1 _5106_/D sky130_fd_sc_hd__clkbuf_1
X_3631_ _3623_/A _3625_/Y _3630_/X vssd1 vssd1 vccd1 vccd1 _3631_/Y sky130_fd_sc_hd__a21oi_1
X_3562_ _3563_/A _3563_/B vssd1 vssd1 vccd1 vccd1 _3562_/X sky130_fd_sc_hd__or2_1
X_2513_ _2515_/A vssd1 vssd1 vccd1 vccd1 _2513_/Y sky130_fd_sc_hd__inv_2
X_5301_ _5301_/A _2500_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
X_3493_ _3494_/A _3494_/B vssd1 vssd1 vccd1 vccd1 _3493_/Y sky130_fd_sc_hd__nand2_1
X_2444_ _2447_/A vssd1 vssd1 vccd1 vccd1 _2444_/Y sky130_fd_sc_hd__inv_2
X_5232_ _5232_/A _2435_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4114_ _4114_/A _4114_/B vssd1 vssd1 vccd1 vccd1 _4116_/A sky130_fd_sc_hd__nand2_1
X_5094_ _5094_/CLK _5094_/D vssd1 vssd1 vccd1 vccd1 _5094_/Q sky130_fd_sc_hd__dfxtp_1
X_4045_ _4993_/Q _4773_/Q vssd1 vssd1 vccd1 vccd1 _4045_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4947_ _4948_/CLK _4947_/D vssd1 vssd1 vccd1 vccd1 _4947_/Q sky130_fd_sc_hd__dfxtp_1
X_4878_ _5058_/CLK _4878_/D vssd1 vssd1 vccd1 vccd1 _4878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3829_ _3829_/A _3829_/B vssd1 vssd1 vccd1 vccd1 _3829_/X sky130_fd_sc_hd__xor2_1
XFILLER_58_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2993_ _2987_/A _2987_/B _2992_/Y vssd1 vssd1 vccd1 vccd1 _2998_/A sky130_fd_sc_hd__o21ai_1
X_4801_ _5015_/CLK _4801_/D vssd1 vssd1 vccd1 vccd1 _4801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4732_ _4942_/Q _5122_/Q _4732_/S vssd1 vssd1 vccd1 vccd1 _4733_/B sky130_fd_sc_hd__mux2_1
X_4663_ _4663_/A vssd1 vssd1 vccd1 vccd1 _5101_/D sky130_fd_sc_hd__clkbuf_1
X_3614_ _3610_/Y _3604_/X _3616_/B _3618_/C _3564_/A vssd1 vssd1 vccd1 vccd1 _3614_/X
+ sky130_fd_sc_hd__a41o_1
X_4594_ _4628_/A vssd1 vssd1 vccd1 vccd1 _4609_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3545_ _3461_/X _3543_/Y _3544_/X _3503_/X vssd1 vssd1 vccd1 vccd1 _4918_/D sky130_fd_sc_hd__o211a_1
X_5165__72 vssd1 vssd1 vccd1 vccd1 _5165__72/HI _5260_/A sky130_fd_sc_hd__conb_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3476_ _3477_/A _3477_/B vssd1 vssd1 vccd1 vccd1 _3476_/X sky130_fd_sc_hd__or2_1
X_2427_ _2428_/A vssd1 vssd1 vccd1 vccd1 _2427_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5077_ _5077_/CLK _5077_/D vssd1 vssd1 vccd1 vccd1 _5077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4028_ _4016_/B _4025_/X _4026_/X _3943_/A vssd1 vssd1 vccd1 vccd1 _4028_/X sky130_fd_sc_hd__a31o_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3330_ _3329_/Y _3309_/B _3307_/Y vssd1 vssd1 vccd1 vccd1 _3330_/Y sky130_fd_sc_hd__a21oi_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5002_/CLK _5000_/D vssd1 vssd1 vccd1 vccd1 _5000_/Q sky130_fd_sc_hd__dfxtp_1
X_3261_ _3254_/B _3259_/X _3260_/X vssd1 vssd1 vccd1 vccd1 _3261_/Y sky130_fd_sc_hd__a21oi_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3192_ _3192_/A _3192_/B vssd1 vssd1 vccd1 vccd1 _3192_/X sky130_fd_sc_hd__and2_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5203__110 vssd1 vssd1 vccd1 vccd1 _5203__110/HI _5311_/A sky130_fd_sc_hd__conb_1
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2976_ _2976_/A vssd1 vssd1 vccd1 vccd1 _2976_/X sky130_fd_sc_hd__clkbuf_2
X_4715_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4730_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4646_ _4646_/A vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__clkbuf_2
X_4577_ _4628_/A vssd1 vssd1 vccd1 vccd1 _4592_/A sky130_fd_sc_hd__clkbuf_2
X_3528_ _3528_/A _3528_/B vssd1 vssd1 vccd1 vccd1 _3529_/C sky130_fd_sc_hd__nand2_1
X_3459_ _4920_/Q _5088_/Q vssd1 vssd1 vccd1 vccd1 _3466_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2830_ _5021_/Q _4813_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _2831_/B sky130_fd_sc_hd__mux2_1
X_2761_ _2761_/A vssd1 vssd1 vccd1 vccd1 _4793_/D sky130_fd_sc_hd__clkbuf_1
X_2692_ _2696_/A _2692_/B vssd1 vssd1 vccd1 vccd1 _2693_/A sky130_fd_sc_hd__and2_1
X_4500_ _4500_/A vssd1 vssd1 vccd1 vccd1 _5054_/D sky130_fd_sc_hd__clkbuf_1
X_4431_ _4855_/Q _5035_/Q _4438_/S vssd1 vssd1 vccd1 vccd1 _4432_/B sky130_fd_sc_hd__mux2_1
XANTENNA_1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5135__42 vssd1 vssd1 vccd1 vccd1 _5135__42/HI _5230_/A sky130_fd_sc_hd__conb_1
X_4362_ _4826_/Q _4814_/Q vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__or2_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _4902_/Q _5070_/Q vssd1 vssd1 vccd1 vccd1 _3327_/A sky130_fd_sc_hd__xor2_2
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _4291_/X _4292_/Y _4230_/X vssd1 vssd1 vccd1 vccd1 _4293_/X sky130_fd_sc_hd__a21o_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3176_/X _3242_/Y _3243_/X _3209_/X vssd1 vssd1 vccd1 vccd1 _4880_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3175_ _3175_/A _3936_/A vssd1 vssd1 vccd1 vccd1 _3182_/A sky130_fd_sc_hd__or2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2959_ _2967_/A _2965_/B _2959_/C vssd1 vssd1 vccd1 vccd1 _4844_/D sky130_fd_sc_hd__nor3_1
XFILLER_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4629_ _4912_/Q _5092_/Q _4629_/S vssd1 vssd1 vccd1 vccd1 _4630_/B sky130_fd_sc_hd__mux2_1
XFILLER_1_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4980_ _4989_/CLK _4980_/D vssd1 vssd1 vccd1 vccd1 _4980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3931_ _4318_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _4021_/B sky130_fd_sc_hd__nor2_2
X_3862_ _4971_/Q _4751_/Q vssd1 vssd1 vccd1 vccd1 _3863_/B sky130_fd_sc_hd__and2_1
X_2813_ _2821_/A _2813_/B vssd1 vssd1 vccd1 vccd1 _2814_/A sky130_fd_sc_hd__and2_1
X_3793_ _3789_/A _3788_/B _3786_/Y vssd1 vssd1 vccd1 vccd1 _3795_/B sky130_fd_sc_hd__a21oi_1
X_2744_ _2744_/A vssd1 vssd1 vccd1 vccd1 _4788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2675_ _2679_/A _2675_/B vssd1 vssd1 vccd1 vccd1 _2676_/A sky130_fd_sc_hd__and2_1
X_4414_ _4850_/Q _5030_/Q _4421_/S vssd1 vssd1 vccd1 vccd1 _4415_/B sky130_fd_sc_hd__mux2_1
X_4345_ _4824_/Q _4812_/Q vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__and2_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4276_ _5022_/Q _4802_/Q vssd1 vssd1 vccd1 vccd1 _4276_/Y sky130_fd_sc_hd__nand2_1
X_3227_ _4891_/Q _5059_/Q vssd1 vssd1 vccd1 vccd1 _3236_/C sky130_fd_sc_hd__or2_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3158_ _3158_/A _3158_/B vssd1 vssd1 vccd1 vccd1 _3160_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3089_ _3083_/A _3083_/B _3088_/Y vssd1 vssd1 vccd1 vccd1 _3094_/A sky130_fd_sc_hd__o21ai_2
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4983_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2460_ input1/X vssd1 vssd1 vccd1 vccd1 _2485_/A sky130_fd_sc_hd__buf_2
X_4130_ _4136_/A vssd1 vssd1 vccd1 vccd1 _4130_/X sky130_fd_sc_hd__clkbuf_2
X_4061_ _4996_/Q _4776_/Q vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__and2_1
XFILLER_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3012_ _2998_/A _2998_/B _3003_/Y _3011_/X vssd1 vssd1 vccd1 vccd1 _3013_/B sky130_fd_sc_hd__a31o_1
XFILLER_36_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _4972_/CLK _4963_/D vssd1 vssd1 vccd1 vccd1 _4963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3914_ _4977_/Q _4757_/Q vssd1 vssd1 vccd1 vccd1 _3915_/B sky130_fd_sc_hd__nand2_1
X_4894_ _5099_/CLK _4894_/D vssd1 vssd1 vccd1 vccd1 _4894_/Q sky130_fd_sc_hd__dfxtp_1
X_3845_ _4969_/Q _4749_/Q vssd1 vssd1 vccd1 vccd1 _3847_/B sky130_fd_sc_hd__xnor2_1
XFILLER_32_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3776_ _4960_/Q _4740_/Q vssd1 vssd1 vccd1 vccd1 _3777_/B sky130_fd_sc_hd__nor2_1
X_2727_ _4992_/Q _4784_/Q _2727_/S vssd1 vssd1 vccd1 vccd1 _2728_/B sky130_fd_sc_hd__mux2_1
X_2658_ _2662_/A _2658_/B vssd1 vssd1 vccd1 vccd1 _2659_/A sky130_fd_sc_hd__and2_1
X_2589_ _2589_/A vssd1 vssd1 vccd1 vccd1 _4744_/D sky130_fd_sc_hd__clkbuf_1
X_4328_ _5017_/Q _4315_/X _4327_/X _4321_/X vssd1 vssd1 vccd1 vccd1 _5017_/D sky130_fd_sc_hd__o211a_1
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4259_ _4306_/B vssd1 vssd1 vccd1 vccd1 _4259_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3630_ _3628_/Y _3630_/B vssd1 vssd1 vccd1 vccd1 _3630_/X sky130_fd_sc_hd__and2b_1
X_3561_ _4933_/Q _5101_/Q vssd1 vssd1 vccd1 vccd1 _3563_/B sky130_fd_sc_hd__xnor2_1
X_2512_ _2515_/A vssd1 vssd1 vccd1 vccd1 _2512_/Y sky130_fd_sc_hd__inv_2
X_5300_ _5300_/A _2499_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3492_ _3477_/A _3477_/B _3483_/Y _3491_/X vssd1 vssd1 vccd1 vccd1 _3494_/B sky130_fd_sc_hd__a31o_1
X_5231_ _5231_/A _2434_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
X_2443_ _2447_/A vssd1 vssd1 vccd1 vccd1 _2443_/Y sky130_fd_sc_hd__inv_2
X_5093_ _5106_/CLK _5093_/D vssd1 vssd1 vccd1 vccd1 _5093_/Q sky130_fd_sc_hd__dfxtp_1
X_4113_ _5002_/Q _4782_/Q vssd1 vssd1 vccd1 vccd1 _4114_/B sky130_fd_sc_hd__nand2_1
X_4044_ _4981_/Q _4034_/X _4043_/Y _4023_/X vssd1 vssd1 vccd1 vccd1 _4981_/D sky130_fd_sc_hd__o211a_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4946_ _4948_/CLK _4946_/D vssd1 vssd1 vccd1 vccd1 _4946_/Q sky130_fd_sc_hd__dfxtp_1
X_4877_ _5058_/CLK _4877_/D vssd1 vssd1 vccd1 vccd1 _4877_/Q sky130_fd_sc_hd__dfxtp_1
X_3828_ _3814_/A _3816_/Y _3821_/B _3819_/Y vssd1 vssd1 vccd1 vccd1 _3829_/B sky130_fd_sc_hd__a31o_1
X_3759_ _4957_/Q _4737_/Q vssd1 vssd1 vccd1 vccd1 _3759_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4800_ _5010_/CLK _4800_/D vssd1 vssd1 vccd1 vccd1 _4800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2992_ _4861_/Q _5029_/Q vssd1 vssd1 vccd1 vccd1 _2992_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4731_ _4731_/A vssd1 vssd1 vccd1 vccd1 _5121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4662_ _4662_/A _4662_/B vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__and2_1
X_3613_ _3610_/Y _3604_/X _3616_/B _3618_/C vssd1 vssd1 vccd1 vccd1 _3613_/Y sky130_fd_sc_hd__a22oi_1
X_4593_ _4593_/A vssd1 vssd1 vccd1 vccd1 _5081_/D sky130_fd_sc_hd__clkbuf_1
X_3544_ _4918_/Q _3544_/B vssd1 vssd1 vccd1 vccd1 _3544_/X sky130_fd_sc_hd__or2_1
X_3475_ _3475_/A _3475_/B vssd1 vssd1 vccd1 vccd1 _3477_/B sky130_fd_sc_hd__and2_1
X_2426_ _2428_/A vssd1 vssd1 vccd1 vccd1 _2426_/Y sky130_fd_sc_hd__inv_2
X_5180__87 vssd1 vssd1 vccd1 vccd1 _5180__87/HI _5288_/A sky130_fd_sc_hd__conb_1
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5076_ _5077_/CLK _5076_/D vssd1 vssd1 vccd1 vccd1 _5076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4027_ _4016_/B _4025_/X _4026_/X vssd1 vssd1 vccd1 vccd1 _4027_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4929_ _5121_/CLK _4929_/D vssd1 vssd1 vccd1 vccd1 _4929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _4895_/Q _5063_/Q vssd1 vssd1 vccd1 vccd1 _3260_/X sky130_fd_sc_hd__xor2_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3191_/A _3191_/B vssd1 vssd1 vccd1 vccd1 _3192_/B sky130_fd_sc_hd__nand2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2975_ _3062_/B vssd1 vssd1 vccd1 vccd1 _2976_/A sky130_fd_sc_hd__buf_2
X_4714_ _4714_/A vssd1 vssd1 vccd1 vccd1 _5116_/D sky130_fd_sc_hd__clkbuf_1
X_4645_ _4645_/A vssd1 vssd1 vccd1 vccd1 _5096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4576_ _4576_/A vssd1 vssd1 vccd1 vccd1 _5076_/D sky130_fd_sc_hd__clkbuf_1
X_3527_ _4928_/Q _5096_/Q vssd1 vssd1 vccd1 vccd1 _3528_/B sky130_fd_sc_hd__or2_1
X_3458_ _4920_/Q _5088_/Q vssd1 vssd1 vccd1 vccd1 _3458_/X sky130_fd_sc_hd__or2_1
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3389_ _3381_/A _3383_/Y _3388_/Y vssd1 vssd1 vccd1 vccd1 _3389_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ _5087_/CLK _5059_/D vssd1 vssd1 vccd1 vccd1 _5059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5077_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2760_ _2767_/A _2760_/B vssd1 vssd1 vccd1 vccd1 _2761_/A sky130_fd_sc_hd__and2_1
X_2691_ _4982_/Q _4774_/Q _2691_/S vssd1 vssd1 vccd1 vccd1 _2692_/B sky130_fd_sc_hd__mux2_1
X_4430_ _4430_/A vssd1 vssd1 vccd1 vccd1 _5034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4361_ _4361_/A vssd1 vssd1 vccd1 vccd1 _4367_/A sky130_fd_sc_hd__clkbuf_2
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _4889_/Q _3277_/A _3310_/Y _3311_/X _3230_/X vssd1 vssd1 vccd1 vccd1 _4889_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _4292_/A _4292_/B vssd1 vssd1 vccd1 vccd1 _4292_/Y sky130_fd_sc_hd__nand2_2
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _4880_/Q _3257_/B vssd1 vssd1 vccd1 vccd1 _3243_/X sky130_fd_sc_hd__or2_1
X_5150__57 vssd1 vssd1 vccd1 vccd1 _5150__57/HI _5245_/A sky130_fd_sc_hd__conb_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3174_ _4884_/Q _5052_/Q vssd1 vssd1 vccd1 vccd1 _3181_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2958_ _4844_/Q _2958_/B vssd1 vssd1 vccd1 vccd1 _2959_/C sky130_fd_sc_hd__and2b_1
X_4628_ _4628_/A vssd1 vssd1 vccd1 vccd1 _4644_/A sky130_fd_sc_hd__clkbuf_2
X_2889_ _2889_/A vssd1 vssd1 vccd1 vccd1 _2889_/X sky130_fd_sc_hd__clkbuf_2
X_4559_ _4646_/A vssd1 vssd1 vccd1 vccd1 _4628_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _4967_/Q _3878_/X _3928_/X _3929_/Y _3866_/X vssd1 vssd1 vccd1 vccd1 _4967_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_16_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3861_ _4971_/Q _4751_/Q vssd1 vssd1 vccd1 vccd1 _3863_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2812_ _5016_/Q _4808_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _2813_/B sky130_fd_sc_hd__mux2_1
X_3792_ _4962_/Q _4742_/Q vssd1 vssd1 vccd1 vccd1 _3805_/A sky130_fd_sc_hd__xor2_1
X_2743_ _2750_/A _2743_/B vssd1 vssd1 vccd1 vccd1 _2744_/A sky130_fd_sc_hd__and2_1
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2674_ _4977_/Q _4769_/Q _2674_/S vssd1 vssd1 vccd1 vccd1 _2675_/B sky130_fd_sc_hd__mux2_1
X_4413_ _4413_/A vssd1 vssd1 vccd1 vccd1 _5029_/D sky130_fd_sc_hd__clkbuf_1
X_4344_ _5019_/Q _4315_/X _4342_/Y _4343_/X _4281_/X vssd1 vssd1 vccd1 vccd1 _5019_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4275_ _5010_/Q _4220_/X _4274_/X _4232_/X vssd1 vssd1 vccd1 vccd1 _5010_/D sky130_fd_sc_hd__o211a_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _4891_/Q _5059_/Q vssd1 vssd1 vccd1 vccd1 _3232_/C sky130_fd_sc_hd__nand2_1
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3157_ _4882_/Q _5050_/Q vssd1 vssd1 vccd1 vccd1 _3158_/B sky130_fd_sc_hd__nand2_1
X_3088_ _4873_/Q _5041_/Q vssd1 vssd1 vccd1 vccd1 _3088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4060_ _4983_/Q _4034_/X _4058_/Y _4059_/X _3962_/X vssd1 vssd1 vccd1 vccd1 _4983_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3011_ _4862_/Q _5030_/Q _3010_/X _3003_/B vssd1 vssd1 vccd1 vccd1 _3011_/X sky130_fd_sc_hd__a31o_1
XFILLER_76_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4962_ _4964_/CLK _4962_/D vssd1 vssd1 vccd1 vccd1 _4962_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3913_ _4977_/Q _4757_/Q vssd1 vssd1 vccd1 vccd1 _3913_/Y sky130_fd_sc_hd__nor2_1
X_4893_ _5087_/CLK _4893_/D vssd1 vssd1 vccd1 vccd1 _4893_/Q sky130_fd_sc_hd__dfxtp_1
X_3844_ _4956_/Q _3838_/X _3843_/X _3797_/X vssd1 vssd1 vccd1 vccd1 _4956_/D sky130_fd_sc_hd__o211a_1
X_3775_ _4960_/Q _4740_/Q vssd1 vssd1 vccd1 vccd1 _3777_/A sky130_fd_sc_hd__and2_1
X_2726_ _2726_/A vssd1 vssd1 vccd1 vccd1 _4783_/D sky130_fd_sc_hd__clkbuf_1
X_2657_ _4972_/Q _4764_/Q _2657_/S vssd1 vssd1 vccd1 vccd1 _2658_/B sky130_fd_sc_hd__mux2_1
X_2588_ _2592_/A _2588_/B vssd1 vssd1 vccd1 vccd1 _2589_/A sky130_fd_sc_hd__and2_1
X_4327_ _4324_/X _4325_/Y _4326_/X vssd1 vssd1 vccd1 vccd1 _4327_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4258_ _4224_/X _4256_/X _4257_/X _4232_/X vssd1 vssd1 vccd1 vccd1 _5008_/D sky130_fd_sc_hd__o211a_1
X_3209_ _4733_/A vssd1 vssd1 vccd1 vccd1 _3209_/X sky130_fd_sc_hd__clkbuf_2
X_4189_ _4189_/A _4189_/B _4191_/C vssd1 vssd1 vccd1 vccd1 _4190_/C sky130_fd_sc_hd__and3_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5186__93 vssd1 vssd1 vccd1 vccd1 _5186__93/HI _5294_/A sky130_fd_sc_hd__conb_1
XFILLER_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3560_ _4920_/Q _3554_/X _3559_/X _3503_/X vssd1 vssd1 vccd1 vccd1 _4920_/D sky130_fd_sc_hd__o211a_1
X_2511_ _2515_/A vssd1 vssd1 vccd1 vccd1 _2511_/Y sky130_fd_sc_hd__inv_2
X_5230_ _5230_/A _2433_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
X_3491_ _4922_/Q _5090_/Q _3490_/X _3483_/B vssd1 vssd1 vccd1 vccd1 _3491_/X sky130_fd_sc_hd__a31o_1
X_2442_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2447_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5092_ _5094_/CLK _5092_/D vssd1 vssd1 vccd1 vccd1 _5092_/Q sky130_fd_sc_hd__dfxtp_1
X_4112_ _5002_/Q _4782_/Q vssd1 vssd1 vccd1 vccd1 _4114_/A sky130_fd_sc_hd__or2_1
X_4043_ _4043_/A _4043_/B vssd1 vssd1 vccd1 vccd1 _4043_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4945_ _5114_/CLK _4945_/D vssd1 vssd1 vccd1 vccd1 _4945_/Q sky130_fd_sc_hd__dfxtp_1
X_4876_ _5058_/CLK _4876_/D vssd1 vssd1 vccd1 vccd1 _4876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3827_ _3827_/A _3827_/B vssd1 vssd1 vccd1 vccd1 _3829_/A sky130_fd_sc_hd__or2_1
X_3758_ _4946_/Q vssd1 vssd1 vccd1 vccd1 _3758_/Y sky130_fd_sc_hd__inv_2
X_2709_ _4987_/Q vssd1 vssd1 vccd1 vccd1 _3992_/A sky130_fd_sc_hd__clkbuf_2
X_3689_ _3712_/A _3689_/B vssd1 vssd1 vccd1 vccd1 _3689_/X sky130_fd_sc_hd__xor2_1
XFILLER_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2991_ _4850_/Q vssd1 vssd1 vccd1 vccd1 _2991_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4730_ _4730_/A _4730_/B vssd1 vssd1 vccd1 vccd1 _4731_/A sky130_fd_sc_hd__and2_1
X_4661_ _4921_/Q _5101_/Q _4665_/S vssd1 vssd1 vccd1 vccd1 _4662_/B sky130_fd_sc_hd__mux2_1
X_3612_ _4939_/Q _5107_/Q vssd1 vssd1 vccd1 vccd1 _3618_/C sky130_fd_sc_hd__or2_1
X_4592_ _4592_/A _4592_/B vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__and2_1
X_3543_ _3546_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3543_/Y sky130_fd_sc_hd__xnor2_1
X_3474_ _4922_/Q _5090_/Q vssd1 vssd1 vccd1 vccd1 _3475_/B sky130_fd_sc_hd__or2_1
X_2425_ _2428_/A vssd1 vssd1 vccd1 vccd1 _2425_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5075_ _5099_/CLK _5075_/D vssd1 vssd1 vccd1 vccd1 _5075_/Q sky130_fd_sc_hd__dfxtp_1
X_4026_ _4991_/Q _4771_/Q vssd1 vssd1 vccd1 vccd1 _4026_/X sky130_fd_sc_hd__xor2_1
X_4928_ _5107_/CLK _4928_/D vssd1 vssd1 vccd1 vccd1 _4928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _5050_/CLK _4859_/D vssd1 vssd1 vccd1 vccd1 _4859_/Q sky130_fd_sc_hd__dfxtp_1
X_5156__63 vssd1 vssd1 vccd1 vccd1 _5156__63/HI _5251_/A sky130_fd_sc_hd__conb_1
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3190_ _3191_/A _3191_/B vssd1 vssd1 vccd1 vccd1 _3192_/A sky130_fd_sc_hd__or2_1
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2974_ _3175_/A _4125_/A vssd1 vssd1 vccd1 vccd1 _3062_/B sky130_fd_sc_hd__nor2_2
XFILLER_34_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4713_ _4713_/A _4713_/B vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5015_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4644_ _4644_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _4645_/A sky130_fd_sc_hd__and2_1
X_4575_ _4575_/A _4575_/B vssd1 vssd1 vccd1 vccd1 _4576_/A sky130_fd_sc_hd__and2_1
X_3526_ _4928_/Q _5096_/Q vssd1 vssd1 vccd1 vccd1 _3528_/A sky130_fd_sc_hd__nand2_1
X_3457_ _3457_/A vssd1 vssd1 vccd1 vccd1 _3457_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3388_ _3388_/A _3388_/B vssd1 vssd1 vccd1 vccd1 _3388_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5058_ _5058_/CLK _5058_/D vssd1 vssd1 vccd1 vccd1 _5058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4009_ _4989_/Q _4769_/Q vssd1 vssd1 vccd1 vccd1 _4010_/B sky130_fd_sc_hd__and2_1
XFILLER_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2690_ _2690_/A vssd1 vssd1 vccd1 vccd1 _4773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4360_ _4319_/X _4358_/Y _4359_/X _4321_/X vssd1 vssd1 vccd1 vccd1 _5021_/D sky130_fd_sc_hd__o211a_1
X_3311_ _3310_/A _3328_/B _3288_/X vssd1 vssd1 vccd1 vccd1 _3311_/X sky130_fd_sc_hd__a21o_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _4292_/A _4292_/B vssd1 vssd1 vccd1 vccd1 _4291_/X sky130_fd_sc_hd__or2_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3242_/A _3245_/A vssd1 vssd1 vccd1 vccd1 _3242_/Y sky130_fd_sc_hd__xnor2_1
X_3173_ _4884_/Q _5052_/Q vssd1 vssd1 vccd1 vccd1 _3173_/X sky130_fd_sc_hd__or2_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2957_ _5285_/A vssd1 vssd1 vccd1 vccd1 _2967_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_41_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2888_ _2886_/X input9/X _2887_/X vssd1 vssd1 vccd1 vccd1 _2888_/X sky130_fd_sc_hd__o21a_1
X_4627_ _4627_/A vssd1 vssd1 vccd1 vccd1 _5091_/D sky130_fd_sc_hd__clkbuf_1
X_4558_ _4558_/A vssd1 vssd1 vccd1 vccd1 _5071_/D sky130_fd_sc_hd__clkbuf_1
X_5126__33 vssd1 vssd1 vccd1 vccd1 _5126__33/HI _5221_/A sky130_fd_sc_hd__conb_1
X_3509_ _3507_/X _3508_/Y _3467_/X vssd1 vssd1 vccd1 vccd1 _3509_/X sky130_fd_sc_hd__a21o_1
X_4489_ _4489_/A vssd1 vssd1 vccd1 vccd1 _5051_/D sky130_fd_sc_hd__clkbuf_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _3851_/Y _3842_/X _3859_/Y _3479_/X vssd1 vssd1 vccd1 vccd1 _4958_/D sky130_fd_sc_hd__a211oi_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2811_ _2811_/A vssd1 vssd1 vccd1 vccd1 _4807_/D sky130_fd_sc_hd__clkbuf_1
X_3791_ _4949_/Q _3784_/X _3789_/Y _3790_/X _3773_/X vssd1 vssd1 vccd1 vccd1 _4949_/D
+ sky130_fd_sc_hd__o221a_1
X_2742_ _4996_/Q _4788_/Q _2745_/S vssd1 vssd1 vccd1 vccd1 _2743_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2673_ _2673_/A vssd1 vssd1 vccd1 vccd1 _4768_/D sky130_fd_sc_hd__clkbuf_1
X_4412_ _4418_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__and2_1
X_4343_ _4333_/A _4336_/B _4341_/Y _4326_/X vssd1 vssd1 vccd1 vccd1 _4343_/X sky130_fd_sc_hd__a31o_1
X_4274_ _4270_/X _4273_/X _4230_/X vssd1 vssd1 vccd1 vccd1 _4274_/X sky130_fd_sc_hd__a21o_1
X_3225_ _3225_/A _3225_/B vssd1 vssd1 vccd1 vccd1 _3225_/X sky130_fd_sc_hd__or2_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3156_ _4882_/Q _5050_/Q vssd1 vssd1 vccd1 vccd1 _3158_/A sky130_fd_sc_hd__or2_1
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3087_ _4862_/Q vssd1 vssd1 vccd1 vccd1 _3087_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _3992_/A _4767_/Q vssd1 vssd1 vccd1 vccd1 _3996_/C sky130_fd_sc_hd__nor2_1
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4966_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3010_ _4863_/Q _5031_/Q vssd1 vssd1 vccd1 vccd1 _3010_/X sky130_fd_sc_hd__or2_1
X_4961_ _4964_/CLK _4961_/D vssd1 vssd1 vccd1 vccd1 _4961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3912_ _4964_/Q _3838_/X _3911_/X _3876_/X vssd1 vssd1 vccd1 vccd1 _4964_/D sky130_fd_sc_hd__o211a_1
X_4892_ _5087_/CLK _4892_/D vssd1 vssd1 vccd1 vccd1 _4892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3843_ _3839_/X _3847_/A _3842_/X vssd1 vssd1 vccd1 vccd1 _3843_/X sky130_fd_sc_hd__a21o_1
X_3774_ _4947_/Q _3745_/X _3771_/Y _3772_/X _3773_/X vssd1 vssd1 vccd1 vccd1 _4947_/D
+ sky130_fd_sc_hd__o221a_1
X_2725_ _2733_/A _2725_/B vssd1 vssd1 vccd1 vccd1 _2726_/A sky130_fd_sc_hd__and2_1
X_2656_ _2656_/A vssd1 vssd1 vccd1 vccd1 _4763_/D sky130_fd_sc_hd__clkbuf_1
X_2587_ _4952_/Q _4744_/Q _2587_/S vssd1 vssd1 vccd1 vccd1 _2588_/B sky130_fd_sc_hd__mux2_1
X_4326_ _4326_/A vssd1 vssd1 vccd1 vccd1 _4326_/X sky130_fd_sc_hd__clkbuf_2
X_4257_ _5008_/Q _4306_/B vssd1 vssd1 vccd1 vccd1 _4257_/X sky130_fd_sc_hd__or2_1
X_4188_ _4999_/Q _4165_/X _4185_/Y _4186_/X _4187_/X vssd1 vssd1 vccd1 vccd1 _4999_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3208_ _4876_/Q _3257_/B vssd1 vssd1 vccd1 vccd1 _3208_/X sky130_fd_sc_hd__or2_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3139_ _4878_/Q _5046_/Q _3139_/C vssd1 vssd1 vccd1 vccd1 _3139_/X sky130_fd_sc_hd__and3_1
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2510_ _2516_/A vssd1 vssd1 vccd1 vccd1 _2515_/A sky130_fd_sc_hd__buf_12
X_3490_ _4923_/Q _5091_/Q vssd1 vssd1 vccd1 vccd1 _3490_/X sky130_fd_sc_hd__or2_1
X_2441_ _2441_/A vssd1 vssd1 vccd1 vccd1 _2441_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4111_ _4989_/Q _4043_/A _4109_/Y _4110_/X _4076_/X vssd1 vssd1 vccd1 vccd1 _4989_/D
+ sky130_fd_sc_hd__o221a_1
X_5091_ _5091_/CLK _5091_/D vssd1 vssd1 vccd1 vccd1 _5091_/Q sky130_fd_sc_hd__dfxtp_1
X_4042_ _4042_/A _4042_/B vssd1 vssd1 vccd1 vccd1 _4043_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4944_ _5114_/CLK _4944_/D vssd1 vssd1 vccd1 vccd1 _4944_/Q sky130_fd_sc_hd__dfxtp_1
X_4875_ _5066_/CLK _4875_/D vssd1 vssd1 vccd1 vccd1 _4875_/Q sky130_fd_sc_hd__dfxtp_1
X_3826_ _4966_/Q _4746_/Q vssd1 vssd1 vccd1 vccd1 _3827_/B sky130_fd_sc_hd__and2_1
X_3757_ _4945_/Q _3745_/X _3756_/X _3724_/X vssd1 vssd1 vccd1 vccd1 _4945_/D sky130_fd_sc_hd__o211a_1
X_2708_ _2708_/A vssd1 vssd1 vccd1 vccd1 _4778_/D sky130_fd_sc_hd__clkbuf_1
X_3688_ _3673_/A _3673_/B _3678_/Y _3687_/X vssd1 vssd1 vccd1 vccd1 _3689_/B sky130_fd_sc_hd__a31o_1
X_2639_ _4967_/Q _4759_/Q _2639_/S vssd1 vssd1 vccd1 vccd1 _2640_/B sky130_fd_sc_hd__mux2_1
X_4309_ _5027_/Q _4807_/Q vssd1 vssd1 vccd1 vccd1 _4309_/Y sky130_fd_sc_hd__xnor2_1
X_5289_ _5289_/A _2484_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
XFILLER_59_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2990_ _4849_/Q _2976_/X _2989_/X _2983_/X vssd1 vssd1 vccd1 vccd1 _4849_/D sky130_fd_sc_hd__o211a_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4660_/A vssd1 vssd1 vccd1 vccd1 _5100_/D sky130_fd_sc_hd__clkbuf_1
X_3611_ _4939_/Q _5107_/Q vssd1 vssd1 vccd1 vccd1 _3616_/B sky130_fd_sc_hd__nand2_1
X_4591_ _4901_/Q _5081_/Q _4595_/S vssd1 vssd1 vccd1 vccd1 _4592_/B sky130_fd_sc_hd__mux2_1
X_3542_ _3528_/A _3530_/X _3535_/B _3533_/Y vssd1 vssd1 vccd1 vccd1 _3543_/B sky130_fd_sc_hd__a31o_1
X_3473_ _4922_/Q _5090_/Q vssd1 vssd1 vccd1 vccd1 _3475_/A sky130_fd_sc_hd__nand2_1
X_2424_ _2428_/A vssd1 vssd1 vccd1 vccd1 _2424_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5074_ _5098_/CLK _5074_/D vssd1 vssd1 vccd1 vccd1 _5074_/Q sky130_fd_sc_hd__dfxtp_1
X_4025_ _4005_/X _4018_/Y _4020_/A _4010_/A vssd1 vssd1 vccd1 vccd1 _4025_/X sky130_fd_sc_hd__a211o_1
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4927_ _5106_/CLK _4927_/D vssd1 vssd1 vccd1 vccd1 _4927_/Q sky130_fd_sc_hd__dfxtp_1
X_4858_ _5040_/CLK _4858_/D vssd1 vssd1 vccd1 vccd1 _4858_/Q sky130_fd_sc_hd__dfxtp_1
X_3809_ _4963_/Q _4743_/Q _4742_/Q _4962_/Q vssd1 vssd1 vccd1 vccd1 _3809_/X sky130_fd_sc_hd__a22o_1
X_4789_ _4999_/CLK _4789_/D vssd1 vssd1 vccd1 vccd1 _4789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5171__78 vssd1 vssd1 vccd1 vccd1 _5171__78/HI _5266_/A sky130_fd_sc_hd__conb_1
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2973_ _4129_/A vssd1 vssd1 vccd1 vccd1 _4125_/A sky130_fd_sc_hd__clkbuf_4
X_4712_ _4936_/Q _5116_/Q _4716_/S vssd1 vssd1 vccd1 vccd1 _4713_/B sky130_fd_sc_hd__mux2_1
X_4643_ _4916_/Q _5096_/Q _4648_/S vssd1 vssd1 vccd1 vccd1 _4644_/B sky130_fd_sc_hd__mux2_1
X_5210__117 vssd1 vssd1 vccd1 vccd1 _5210__117/HI _5318_/A sky130_fd_sc_hd__conb_1
X_4574_ _4896_/Q _5076_/Q _4578_/S vssd1 vssd1 vccd1 vccd1 _4575_/B sky130_fd_sc_hd__mux2_1
X_3525_ _3494_/A _3494_/B _3522_/Y _3524_/Y _3521_/B vssd1 vssd1 vccd1 vccd1 _3529_/B
+ sky130_fd_sc_hd__a311oi_2
X_3456_ _3544_/B vssd1 vssd1 vccd1 vccd1 _3457_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3387_ _4911_/Q _5079_/Q vssd1 vssd1 vccd1 vccd1 _3388_/B sky130_fd_sc_hd__and2_1
XFILLER_84_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5057_ _5058_/CLK _5057_/D vssd1 vssd1 vccd1 vccd1 _5057_/Q sky130_fd_sc_hd__dfxtp_1
X_4008_ _4989_/Q _4769_/Q vssd1 vssd1 vccd1 vccd1 _4010_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5066_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3310_ _3310_/A _3328_/B vssd1 vssd1 vccd1 vccd1 _3310_/Y sky130_fd_sc_hd__nor2_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ _4290_/A _4290_/B vssd1 vssd1 vccd1 vccd1 _4292_/B sky130_fd_sc_hd__and2_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1 _3245_/A sky130_fd_sc_hd__nand2_1
X_3172_ _3223_/A vssd1 vssd1 vccd1 vccd1 _3172_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ _2956_/A vssd1 vssd1 vccd1 vccd1 _4843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2887_ _2905_/A vssd1 vssd1 vccd1 vccd1 _2887_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4626_ _4626_/A _4626_/B vssd1 vssd1 vccd1 vccd1 _4627_/A sky130_fd_sc_hd__and2_1
X_4557_ _4557_/A _4557_/B vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__and2_1
X_3508_ _3521_/A _3508_/B vssd1 vssd1 vccd1 vccd1 _3508_/Y sky130_fd_sc_hd__nand2_1
X_4488_ _4488_/A _4488_/B vssd1 vssd1 vccd1 vccd1 _4489_/A sky130_fd_sc_hd__and2_1
X_3439_ _3430_/A _3432_/Y _3438_/X vssd1 vssd1 vccd1 vccd1 _3439_/Y sky130_fd_sc_hd__a21oi_1
X_5141__48 vssd1 vssd1 vccd1 vccd1 _5141__48/HI _5236_/A sky130_fd_sc_hd__conb_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5109_ _5121_/CLK _5109_/D vssd1 vssd1 vccd1 vccd1 _5109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2810_ _2821_/A _2810_/B vssd1 vssd1 vccd1 vccd1 _2811_/A sky130_fd_sc_hd__and2_1
X_3790_ _3789_/A _3806_/B _3755_/X vssd1 vssd1 vccd1 vccd1 _3790_/X sky130_fd_sc_hd__a21o_1
X_2741_ _2741_/A vssd1 vssd1 vccd1 vccd1 _4787_/D sky130_fd_sc_hd__clkbuf_1
X_2672_ _2679_/A _2672_/B vssd1 vssd1 vccd1 vccd1 _2673_/A sky130_fd_sc_hd__and2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4411_ _4849_/Q _5029_/Q _4421_/S vssd1 vssd1 vccd1 vccd1 _4412_/B sky130_fd_sc_hd__mux2_1
X_4342_ _4333_/A _4336_/B _4341_/Y vssd1 vssd1 vccd1 vccd1 _4342_/Y sky130_fd_sc_hd__a21oi_1
X_4273_ _4284_/A _4256_/B _4263_/A _4283_/A _4272_/Y vssd1 vssd1 vccd1 vccd1 _4273_/X
+ sky130_fd_sc_hd__a311o_1
X_3224_ _4878_/Q _3172_/X _3223_/Y _3209_/X vssd1 vssd1 vccd1 vccd1 _4878_/D sky130_fd_sc_hd__o211a_1
.ends

